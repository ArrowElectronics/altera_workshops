-- top.vhd

-- Generated using ACDS version 24.2 40

library IEEE;
library altera_mult_add_1921;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity top_answer is
	port (
		dataa : in  std_logic_vector(15 downto 0)  := (others => '0'); -- dataa_0.dataa_0, Input a of multiplier-adder
		datab : in  std_logic_vector(15 downto 0)  := (others => '0'); -- dataa_0.dataa_0, Input a of multiplier-adder
		denom : in  std_logic_vector(15 downto 0)  := (others => '0'); -- dataa_0.dataa_0, Input a of multiplier-adder
		result  : out std_logic_vector(31 downto 0);                    --  result.result,  Result of the multiplier-adder
		remain : out std_logic_vector(15 downto 0)  ; 
		clock0  : in  std_logic                      := '0';              --  clock0.clk,     Clock input port to the corresponding register. This port can be used by any register in the IP core.
		clock1  : in  std_logic                      := '0'              --  clock1.clk,     Clock input port to the corresponding register. This port can be used by any register in the IP core.		
	
	);

end entity top_answer;

architecture rtl of top_answer is

		component Div32by16 is
		port (
			numer    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- numer
			denom    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- denom
			clock    : in  std_logic                     := 'X';             -- clock
			quotient : out std_logic_vector(31 downto 0);                    -- quotient
			remain   : out std_logic_vector(15 downto 0)                     -- remain
		);
	end component Div32by16;

	component Mult16x16 is
		port (
			dataa  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- dataa
			result : out std_logic_vector(31 downto 0);                    -- result
			datab  : in  std_logic_vector(15 downto 0) := (others => 'X')  -- datab
		);
	end component Mult16x16;

	
	
	signal mult_result    : std_logic_vector(31 downto 0);     
	signal mult_result_r  : std_logic_vector(31 downto 0);     
	signal dataa_r : std_logic_vector(15 downto 0);     -- datab_0.datab_0, Input b of multiplier-adder
	signal datab_r : std_logic_vector(15 downto 0);     -- datab_0.datab_0, Input b of multiplier-adder
	signal dataa_r1 : std_logic_vector(15 downto 0);     -- datab_0.datab_0, Input b of multiplier-adder
	signal datab_r1 : std_logic_vector(15 downto 0);     -- datab_0.datab_0, Input b of multiplier-adder
	signal denom_r : std_logic_vector(15 downto 0)  := (others => '0'); -- dataa_0.dataa_0, Input a of multiplier-adder
	signal result_u : std_logic_vector(31 downto 0);     -- datab_0.datab_0, Input b of multiplier-adder
	signal remain_u : std_logic_vector(15 downto 0)  := (others => '0'); -- dataa_0.dataa_0, Input a of multiplier-adder
	signal denom_r0 : std_logic_vector(15 downto 0);
	signal denom_r1 : std_logic_vector(15 downto 0);
	signal denom_r2 : std_logic_vector(15 downto 0);

	
begin

	CAPTURE_DATA0 : process (clock1)
	begin	
		if rising_edge(clock1) then
			dataa_r <= dataa;
			datab_r <= datab;
		end if;
	end process CAPTURE_DATA0;
	
	CAPTURE_DATA1 : process (clock0)
	begin	
		if rising_edge(clock0) then
			dataa_r1 <= dataa_r;
			datab_r1 <= datab_r;
			denom_r <= denom;
			denom_r0 <= denom_r;
			denom_r1 <= denom_r0;
			denom_r2 <= denom_r1;
		end if;
	end process CAPTURE_DATA1;
	
	CAPTURE_OUT0 : process (clock0)
	begin	
		if rising_edge(clock0) then
			mult_result_r <= mult_result;
			result <= result_u;
			remain <= remain_u;
		end if;
	end process CAPTURE_OUT0;
	
	

	u0 : component Mult16x16
		port map (
			dataa  => dataa_r1,  --  dataa.dataa
			result => mult_result, -- result.result
			datab  => datab_r1   --  datab.datab
		);
	
	u1 : component Div32by16
		port map (
			numer    => mult_result_r,    --  lpm_divide_input.numer
			denom    => denom_r2,    --                  .denom
			clock    => clock0,             -- clock
			quotient => result_u, -- lpm_divide_output.quotient
			remain   => remain_u    --                  .remain
		);
	
	

end architecture rtl; -- of top

----------------------------------------------------------------
-- SPDX-FileCopyrightText: Copyright (C) 2025 Arrow Electronics, Inc. 
-- SPDX-License-Identifier: MIT-0 
----------------------------------------------------------------
--
--Design Name:		SignalTap Lab
--Module Name:		Top module
--Version:			1.0
--Created Date:		18 June 2024
--
--Company:			Arrow Electronics
--Author:			Szabolcs Bondor
--
--Configuration:
--Target Device:	Altera Agilex5 E-Series
--Target Board:	Arrow AXE5-Eagle Board
--Software:			Quartus Prime Pro 24.1
--
--Description:		This lab realizes a simple UART TX interface 
--						without parity bit. For the parallel-serial 
--						conversion it uses a shift register, while the 
--						data is generated by a counter.
--						
--Note:				
--History:			Fue Xiong: Repurposed top level design file for the Arrow AXE5-Eagle Board
--  					Updated IP instance to align with IP variants from Prime Pro
----------------------------------------------------------------


---------------------------[LIBRARY]----------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

---------------------------[ENTITY]-----------------------------

entity uart_tx is
port(	CLK			: in std_logic;
--***** uncomment the next line of code if using local hardware
--		BTN			: in std_logic;
		UART_TX		: out std_logic);
end entity uart_tx;

------------------------[ARCHITECTURE]--------------------------

architecture Behavioral of uart_tx is

signal nINIT_DONE   	: std_logic;
signal iCLK			    : std_logic;
signal iCTRL		    : std_logic := '0';
signal iDATACNT	    	: std_logic_vector(7 downto 0);
signal iDATASHFT	  	: std_logic_vector(0 to 7);

signal clks_per_bit		: integer := 217;
signal clk_cnt       	: integer range 0 to clks_per_bit-1 := 0;
signal baud_out      	: std_logic;

signal BTNn             : std_logic;
signal iDATASHFT_concat : std_logic_vector(0 to 9);

--***** uncomment the next two lines of code if using board farm hardware
--signal jtag_src			: std_logic_vector(0 to 0);
--signal BTN		  		: std_logic;

----------------------------------------------------------------
--                                                            --
--           RESET RELEASE COMPONENT DECLARATION              --
--                  INSERT TEMPLATES BELOW                    --
--                                                            --
----------------------------------------------------------------
	component reset_release is
		port (
			ninit_done : out std_logic   -- reset
		);
	end component reset_release;

----------------------------------------------------------------
--                                                            --
--                 PLL COMPONENT DECLARATION                  --
--                  INSERT TEMPLATES BELOW                    --
--                                                            --
----------------------------------------------------------------
	component PLL is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic         -- clk
		);
	end component PLL;

----------------------------------------------------------------
--                                                            --
--               COUNTER COMPONENT DECLARATION                --
--                  INSERT TEMPLATES BELOW                    --
--                                                            --
----------------------------------------------------------------
	component counter is
		port (
			clock  : in  std_logic                    := 'X';             -- clock
			cnt_en : in  std_logic                    := 'X';             -- cnt_en
			sload  : in  std_logic                    := 'X';             -- sload
			data   : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			q      : out std_logic_vector(7 downto 0)                     -- q
		);
	end component counter;

----------------------------------------------------------------
--                                                            --
--            SHIFT REGISTER COMPONENT DECLARATION            --
--                  INSERT TEMPLATES BELOW                    --
--                                                            --
----------------------------------------------------------------
	component shiftregister is
		port (
			clock    : in  std_logic                    := 'X';             -- clock
			load     : in  std_logic                    := 'X';             -- load
			data     : in  std_logic_vector(9 downto 0) := (others => 'X'); -- data
			sset     : in  std_logic                    := 'X';             -- sset
			shiftout : out std_logic                                        -- shiftout
		);
	end component shiftregister;
	
----------------------------------------------------------------
--                                                            --
--             JTAG SOURCECOMPONENT DECLARATION            	  --
--                  INSERT TEMPLATES BELOW                    --
--                                                            --
----------------------------------------------------------------
--***** uncomment the next five lines of code if using board farm hardware	
--	component jtag_source is
--		port (
--			source : out std_logic_vector(0 downto 0)
--		);
--	end component jtag_source;

begin

   SDM_INIT_DONE : reset_release
   port map (
     ninit_done => nINIT_DONE  -- ninit_done.reset
   );


	clock : PLL
	port map(refclk   => CLK,
	         rst      => nINIT_DONE,
				   outclk_0 => iCLK);
	
	
	datagen : counter
	port map(clock  => baud_out,
				   cnt_en => '1',
				   sload  => '0',				
				   data   => x"56",
				   q      => iDATACNT);
	
	
	serdes : shiftregister
	port map(clock    => baud_out,
				   load     => iCTRL,	
				   data     => iDATASHFT_concat,
				   sset     => BTNn,
				   shiftout => UART_TX);

  BTNn             <= not BTN;
  iDATASHFT_concat <= '0' & iDATASHFT & '1';
				
	load : process(baud_out, BTN)
	variable delay : std_logic_vector(3 downto 0) := x"F";
	begin
		if (BTN = '0') then
			delay := x"F";
			iCTRL <= '0';
		elsif (baud_out = '0' and baud_out'event) then
			if (delay = x"F") then
				iCTRL <= '1';
				delay := x"0";
			else
				iCTRL <= '0';
				delay := delay + 1;
			end if;
		end if;
	end process;

  -- Generate pulse for baudrate
  -- Since the input clock is much faster than the baudrate of the UART interface,
  -- to not over transmit data, count the number of clocks per bit transfer and
  -- generate a pulse to represent the baudrate clock.
  -- Ex. CLK=25Mhz, Baudrate=115200, 25000000/115200=217 clocks per bit
	baud_rate : process (iCLK, nINIT_DONE)
  begin
    if(nINIT_DONE = '1') then
      clk_cnt  <= 0;
      baud_out <= '0';
    elsif(rising_edge(iCLK)) then
      if (clk_cnt = clks_per_bit-1) then
        clk_cnt <= 0;
        baud_out <= not baud_out;
      else
        clk_cnt <= clk_cnt + 1;
      end if;
    end if;
  end process;
  
  
	reverse : process (iDATACNT)
	begin
		for i in iDATACNT'range loop
			iDATASHFT(i) <= iDATACNT(i);
		end loop;
	end process;

--***** uncomment the next five lines of code if using board farm hardware	
--	u4 : jtag_source	
--	port map (
--		source => jtag_src
--	);

--	BTN <= jtag_src(0);
	

	
end architecture Behavioral;

-----------------------------[END]------------------------------

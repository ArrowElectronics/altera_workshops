library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
use work.CNN_Config_Package.all;
use work.CNN_Data_Package.all;

PACKAGE Test_Data_Package is

  type Image_Array_T is array (0 to 127, 0 to 127) of CNN_Values_T (2 downto 0);

  CONSTANT Image_Example : Image_Array_T :=
  (
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (0, 0, 0), (0, 0, 0), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127)),
    ((127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127), (127, 127, 127))
  );
END PACKAGE Test_Data_Package;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
use work.CNN_Config_Package.all;

PACKAGE CNN_Data_Package is
  CONSTANT Layer_1_Columns    : NATURAL := 128;
  CONSTANT Layer_1_Rows       : NATURAL := 128;
  CONSTANT Layer_1_Strides    : NATURAL := 1;
  CONSTANT Layer_1_Activation : Activation_T := relu;
  CONSTANT Layer_1_Padding    : Padding_T := same;
  CONSTANT Layer_1_Values     : NATURAL := 1;
  CONSTANT Layer_1_Filter_X   : NATURAL := 3;
  CONSTANT Layer_1_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_1_Filters    : NATURAL := 12;
  CONSTANT Layer_1_Inputs     : NATURAL := 10;
  CONSTANT Layer_1_Out_Offset : INTEGER := 3;
  CONSTANT Layer_1_Offset     : INTEGER := 0;
  CONSTANT Layer_1 : CNN_Weights_T(0 to Layer_1_Filters-1, 0 to Layer_1_Inputs-1) :=
  (
    (-79, -84, -78, -31, 4, 74, 68, 37, 36, -3),
    (28, 61, 69, 2, 6, -30, -81, -124, -35, -1),
    (-40, -27, 23, -66, 73, -22, 79, 83, 40, 4),
    (-51, -27, -6, -25, -13, 41, -50, 14, -52, 1),
    (87, 5, 68, 29, -54, 94, -50, 27, -35, 1),
    (42, -13, -59, 51, -4, 32, 22, 61, 69, -11),
    (99, 26, -121, -41, 0, -41, -60, -5, -51, -1),
    (-26, 22, -85, -14, -39, -77, 117, 5, -85, 1),
    (67, 4, 72, 81, -1, 100, -28, -41, 41, -9),
    (-78, -45, 74, -88, -11, 86, 41, 27, 5, 3),
    (-41, 74, -64, -50, 56, 64, -82, 40, -104, 1),
    (110, -71, -67, 36, -99, -16, -15, 21, 10, -5)
  );
  ----------------
  CONSTANT Pooling_1_Columns      : NATURAL := 128;
  CONSTANT Pooling_1_Rows         : NATURAL := 128;
  CONSTANT Pooling_1_Values       : NATURAL := 12;
  CONSTANT Pooling_1_Filter_X     : NATURAL := 2;
  CONSTANT Pooling_1_Filter_Y     : NATURAL := 2;
  CONSTANT Pooling_1_Strides      : NATURAL := 2;
  CONSTANT Pooling_1_Padding      : Padding_T := valid;
  ----------------
  CONSTANT Layer_2_Columns    : NATURAL := 64;
  CONSTANT Layer_2_Rows       : NATURAL := 64;
  CONSTANT Layer_2_Strides    : NATURAL := 2;
  CONSTANT Layer_2_Activation : Activation_T := relu;
  CONSTANT Layer_2_Padding    : Padding_T := same;
  CONSTANT Layer_2_Values     : NATURAL := 12;
  CONSTANT Layer_2_Filter_X   : NATURAL := 3;
  CONSTANT Layer_2_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_2_Filters    : NATURAL := 16;
  CONSTANT Layer_2_Inputs     : NATURAL := 109;
  CONSTANT Layer_2_Out_Offset : INTEGER := 3;
  CONSTANT Layer_2_Offset     : INTEGER := 0;
  CONSTANT Layer_2 : CNN_Weights_T(0 to Layer_2_Filters-1, 0 to Layer_2_Inputs-1) :=
  (
    (-26, 38, -17, -50, 21, -18, -9, 1, 13, 6, 10, 12, -31, 45, -11, -28, 39, -12, -5, -10, 11, -4, -2, -3, -33, 51, -15, -44, 34, -18, 7, -5, 1, 7, 1, -1, 33, 30, -6, -15, -25, -21, -13, 20, -20, 17, -20, 29, 47, 36, 16, -21, -24, -28, 19, 12, -8, -4, -32, 14, 14, 15, 4, -3, -21, -6, 25, 14, -5, 2, -5, 8, -9, -24, 0, -41, -7, 34, -30, 0, 14, 4, -24, -15, 7, 6, 10, -32, 1, 23, -48, -10, -5, -2, -27, -13, 27, 10, 23, -14, -6, 12, -6, -4, 0, -6, -25, -19, -2),
    (29, 10, -4, 13, -38, -21, -18, 22, 12, 3, 0, 29, -30, 9, 12, 24, 6, -35, -15, 24, -19, 22, 23, -20, -39, 43, -3, 17, 12, -7, -17, -47, 26, 39, 11, -14, 26, -41, 2, -13, -14, -8, -2, 55, 12, -2, -8, 13, 9, 40, -10, 62, -23, 2, -42, 55, -23, 14, -1, -3, -35, 28, -12, -8, 24, 7, -43, 2, -14, 29, 22, -56, 1, -46, 3, -12, -17, 10, -25, 56, 33, -9, 17, 34, 19, -10, 23, 34, -23, 2, -30, 32, -8, -28, 15, 20, 14, 0, -24, 44, 0, -16, -46, -11, 8, -6, -9, 4, 2),
    (15, 13, 10, -47, 5, -31, -13, 0, -10, 31, -37, 8, 1, -15, 16, -78, -26, -3, 6, 15, 30, 20, -33, 33, -22, 5, 9, -38, -1, 4, -14, 23, 26, 7, -20, 21, 10, 11, 18, -75, -28, -26, 3, -18, 12, 35, -38, 33, 27, 1, 4, -64, 4, -13, 16, -6, -18, 30, -29, 48, 8, 3, 22, -17, -5, -15, -5, -17, 5, 10, -7, 24, -10, -12, -30, -44, -27, -10, 0, -1, -17, 39, -4, 35, -13, 20, 24, -79, 1, 12, 18, 2, -26, 36, -29, 48, 18, 20, 22, -16, 13, 19, 8, -9, 21, 3, -2, 29, -2),
    (9, 1, 27, -1, -20, 21, 17, -9, -19, -1, -5, 25, 13, -1, -19, 24, -26, -20, -3, 37, -13, -23, 31, 29, 8, -2, 14, 25, 12, 3, -15, 49, -29, -7, 19, 22, 26, 60, -3, -8, -3, -31, 11, -27, 14, -15, 22, -3, -12, 10, -18, -1, -2, -8, 21, -19, 10, 12, 43, -1, -11, 12, 20, 17, -6, 15, 6, -15, 14, 6, 8, 7, 20, 36, -4, -24, 11, -29, -20, 4, 3, 2, 34, 8, -31, 0, -31, -17, 13, -22, 7, 5, -7, 10, 12, 10, -27, 25, -4, -10, 1, -31, 12, -33, 30, -24, -3, -10, -1),
    (-22, 31, 16, -24, 24, 26, 37, 18, 11, -15, -10, 30, -40, -6, 10, 5, -3, 14, 40, 2, 8, -22, -8, 31, 3, 14, 7, 13, -6, -29, 17, -17, -10, -7, -30, 30, -1, 21, -8, 13, -24, 5, 29, -10, 14, 4, -15, 30, 20, -2, -24, 11, 6, -23, 32, 20, -31, 21, -26, 28, 27, -17, 6, 0, -11, 0, 21, -36, -21, 16, -37, 22, 7, 21, 12, 1, -25, -22, -8, -14, -16, -6, -23, 12, 17, -29, -14, 1, 5, -11, 4, -19, -34, 21, -36, -14, 8, -19, 3, -6, 6, 29, -44, -5, 31, 34, -10, -18, 4),
    (23, 22, -13, 22, -2, -27, 2, -4, -4, 6, -2, -6, -11, 10, -13, -30, 8, 12, -12, -12, 4, -13, -9, -11, -23, 12, -10, -22, 27, 21, -1, -4, 18, -10, 9, -14, -1, -22, 29, 16, -33, -2, -33, 28, 3, 13, -33, 14, 5, 23, -21, 17, -10, -19, -7, 20, -17, 25, -13, -37, -16, 14, -12, 3, -18, 4, 20, -36, -8, -10, -21, 17, -3, -27, 3, -34, -22, 33, 6, 28, 1, 13, -7, -4, 12, -21, -13, 3, -19, 2, -15, 19, -16, -28, -3, -2, -15, -14, -39, 2, -15, -26, -30, 8, -25, -1, 2, 4, -1),
    (13, 27, 17, -22, -16, -8, 8, -12, -10, -28, -8, -18, -3, -3, 23, -39, -14, 32, -9, 2, 18, -30, 12, -25, 16, 12, -18, -27, 3, 2, -9, -23, 9, -7, 19, 5, -10, -11, -12, -11, 18, 46, -1, -15, -8, -13, 12, -11, 4, 8, 29, -13, 2, 8, -17, -48, 17, -33, -8, -42, 5, -8, 32, 8, 4, 1, -38, -38, -4, -11, 8, -16, -21, -3, 11, 4, 27, 30, -20, -23, 33, -16, 4, -1, -17, -2, 12, -27, 5, 25, -20, -29, 4, -23, 9, -3, -25, 6, 20, -37, -8, -8, -13, 6, 29, -20, -1, -22, -3),
    (-4, 38, 7, -13, 24, 7, -17, -13, 15, -13, 26, -2, 2, -7, 5, -22, -9, -27, 1, 15, -4, 22, -7, 17, -1, -10, 13, -24, 4, -12, 15, 16, -23, -39, 10, -13, 16, -10, -23, 42, -14, 6, -19, 1, -7, 4, -9, -14, 2, 7, -11, 24, -11, -33, -3, -4, -34, 21, -3, -21, 27, -27, -18, -16, -8, -28, 5, 38, 3, -13, -28, 0, 28, 23, 30, 6, -14, -5, -15, 9, 16, 12, -1, -18, 20, -6, 30, 30, -24, 4, 23, -3, -31, 0, -11, -8, 10, -8, 32, 15, -20, -23, -28, 19, -7, -26, 32, 33, 0),
    (-35, -14, 22, -38, 28, -5, -10, -10, 18, 1, 6, -5, -39, -20, 31, -40, 6, 39, -22, 2, -1, 3, 11, 13, -1, -3, 1, -51, 29, 39, 13, 1, 20, 5, 9, 11, -48, -24, -26, 36, 12, -14, 19, -4, 12, -4, 13, 22, -27, -11, 9, 7, 23, 28, 15, 2, 4, -12, 6, -30, -39, -18, -2, -1, 12, 20, -3, -10, -15, 10, 17, -15, -41, -12, -30, -8, 10, 9, 4, 0, 7, 19, 3, 4, -35, -14, 1, 1, 0, 23, 14, 6, 6, -25, 24, 9, -19, -16, -12, 8, -6, 30, 18, 10, -2, -19, 31, -11, 2),
    (-5, 2, 18, -27, 9, 4, 0, -10, 32, -10, -1, -9, -3, 7, 7, -50, -4, -3, 2, -33, 40, 5, 7, -21, -10, -9, -7, -69, -7, 14, -10, -30, 18, 10, 4, -14, -13, 29, -40, -67, -1, 9, 4, -15, -1, 11, 19, -5, -16, 56, -28, -49, 28, -30, -11, -30, 19, -2, 12, -3, -1, 36, -31, -30, 33, -24, -18, -22, 30, -2, -3, -7, 39, 21, 11, 3, -21, 0, 5, 7, -39, -17, -6, 18, 29, 47, -21, -23, -20, 8, -12, 12, -22, 20, 6, 20, 34, 25, -1, 3, 14, -16, 18, 1, -32, -1, -2, 4, -1),
    (-34, -21, 19, -46, -31, 11, -7, -13, 12, 3, -11, 13, -7, -13, 4, -93, 3, -13, 7, -18, 29, 15, -2, 36, -12, -9, 14, 1, -1, 0, -14, -1, -15, 11, -19, 17, -32, -28, 33, -47, 22, 8, 17, -3, 1, -6, -24, 39, -30, -5, 13, -93, -7, 26, 12, 8, 11, 24, 5, 29, -3, 25, 18, -56, 17, 24, -14, 1, -1, 14, -8, 11, -25, -2, 19, -16, 3, -5, 11, 11, 24, -19, -5, 28, -20, 8, 16, -59, -18, -2, -1, -5, 33, 10, -17, 38, 20, 32, 7, -40, 3, 17, -24, -15, 18, 7, -8, 26, -2),
    (1, 36, -11, 41, -20, -9, -22, 23, -33, -2, 16, 10, -1, 41, -29, 14, -10, -36, -27, 27, -13, -13, 8, -8, -29, 13, -18, 11, 7, -28, -29, 20, -5, 0, 10, -50, 12, 40, 28, -18, -16, -4, -12, -6, 18, -5, -18, -10, 0, -6, -1, 18, 9, 2, 0, 43, -1, 9, 5, -12, 0, 34, 17, 29, 11, -10, -35, 26, -23, -9, 10, 8, -21, 19, -10, -15, 30, 35, 3, -6, 5, 13, 11, -10, -2, 11, 28, -16, 15, 31, -9, 38, -10, -18, 0, -17, 0, -32, 9, 14, -5, 35, -20, 23, -14, 0, -7, 3, 0),
    (4, -24, 8, 40, -16, 6, 17, -15, 9, 16, 27, -5, -3, -20, 21, -10, -35, 5, 3, 5, 5, 21, 17, -18, 21, -25, 25, -7, -21, -26, -12, 8, -31, -35, 11, 16, 4, 33, 21, 29, -7, 9, 11, 16, -14, 8, 14, 4, 31, 30, 16, -12, 10, -2, 18, 21, 28, 0, 37, 4, -9, 1, -31, 6, 13, -26, -9, 13, -36, 2, -28, 31, 23, 8, 31, 24, -15, -34, 18, -1, 13, 11, -17, 15, 5, 43, -29, -27, -11, 14, 4, 16, -5, 3, -30, -23, -50, -9, -34, -15, -28, -42, -22, -4, -5, -17, -46, 24, 4),
    (1, -65, 34, -52, 5, 36, -23, -14, -13, 17, -1, -18, 11, -37, 15, -19, 9, -10, 4, -41, -13, -11, -13, -13, -20, -51, 8, -10, 3, 16, 27, -29, -23, 8, -20, 0, 14, -2, 5, -24, -16, 20, 1, -7, -5, -7, -28, -23, -29, -30, 26, -77, -14, 26, -18, -31, 37, 6, 6, 6, -10, -14, 11, -35, -2, -4, 4, -16, 13, -12, -18, 8, -6, -32, 6, -51, 0, 21, 1, -1, 23, 7, -25, 31, 12, -22, -2, -63, 7, 30, -6, -9, -19, -10, -13, -12, 9, -11, 17, -22, 11, 12, -5, -23, 14, -14, -21, -11, -2),
    (-23, -4, -22, 25, -35, 17, 21, -20, -6, 13, 8, 0, -13, 15, 9, 37, 23, -34, 42, 8, -23, 8, -5, -3, 1, -11, -18, -2, 25, 20, 18, -3, -14, -9, 11, 24, 29, -21, 2, 26, -20, 1, 0, -13, -32, -19, -4, 18, -26, -32, 22, 11, -4, 12, -34, -6, -22, -9, -33, -11, -17, 6, -15, -1, -4, -29, -29, -21, -8, -8, 35, 15, -3, 50, 14, 26, 5, -22, 6, -25, 23, -34, 23, 6, -7, 4, 21, 30, 5, -6, 8, 3, 5, 1, -18, -27, -10, -21, -13, -17, -8, 8, 13, -8, 6, 9, -11, 22, -2),
    (6, -23, -2, -2, -13, 28, 1, 2, 13, -11, -37, -14, 21, 7, 16, -5, -18, -9, -4, 9, 5, 2, -20, 4, 1, -28, -3, -4, -26, 11, -10, -6, -7, -31, -27, -16, 4, -29, 18, -41, 1, 39, -2, 27, -9, -24, -18, -12, 25, -7, -10, -3, -23, 16, -30, -5, -12, 11, -7, -5, 16, -46, -5, 4, -20, -7, 12, 32, -16, -6, -28, 3, -22, -35, 20, 10, 25, 7, -18, 21, -8, 30, 5, 28, -11, -35, -8, -31, 26, 2, -25, 26, -4, -8, -3, 27, 26, -32, 0, 20, -23, -7, -10, 9, -27, -11, -16, 2, -2)
  );
  ----------------
  CONSTANT Layer_3_Columns    : NATURAL := 32;
  CONSTANT Layer_3_Rows       : NATURAL := 32;
  CONSTANT Layer_3_Strides    : NATURAL := 2;
  CONSTANT Layer_3_Activation : Activation_T := relu;
  CONSTANT Layer_3_Padding    : Padding_T := same;
  CONSTANT Layer_3_Values     : NATURAL := 16;
  CONSTANT Layer_3_Filter_X   : NATURAL := 3;
  CONSTANT Layer_3_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_3_Filters    : NATURAL := 24;
  CONSTANT Layer_3_Inputs     : NATURAL := 145;
  CONSTANT Layer_3_Out_Offset : INTEGER := 3;
  CONSTANT Layer_3_Offset     : INTEGER := -1;
  CONSTANT Layer_3 : CNN_Weights_T(0 to Layer_3_Filters-1, 0 to Layer_3_Inputs-1) :=
  (
    (-1, 22, 11, -4, 21, 18, -41, -38, 25, 30, -56, 62, 41, -60, -36, 11, -18, 72, -14, -25, -72, -3, -27, 13, -41, -32, -39, 13, 56, -75, -11, 37, 6, 53, 26, 32, -16, -43, -7, -13, 68, 10, 60, 42, -100, 21, -44, -1, -9, 41, -16, 41, -32, 34, -20, 32, 48, 4, 38, 52, 2, 24, 2, 50, 5, 45, -51, -19, -89, -4, -39, 10, -60, -30, -31, 46, -12, -7, 20, 50, -42, 78, 58, 46, 24, -55, -26, -82, 28, 44, -9, -5, -55, -20, -90, -67, -10, 27, 38, -27, -72, 12, -40, 3, 59, -54, -23, 4, -9, -25, -11, 62, -2, 52, -35, -32, -22, 12, 27, -10, -19, -21, 11, 46, 3, 66, -10, 46, 23, 42, 36, 31, -16, 6, 3, -27, -28, 63, -21, -23, -19, -38, -8, -48, -8),
    (30, 48, 8, 36, -14, 62, -21, -13, 49, 40, 2, 66, 17, 31, 63, -58, -10, 44, -32, 10, -33, 86, 53, -30, 28, 75, -26, 49, 17, 9, 32, -27, -18, 100, -19, 62, -43, -21, 61, 31, 55, 38, -24, 82, -29, 23, 38, 17, 2, 1, 1, -86, -22, 107, -23, -25, -27, 9, 7, 3, -65, -23, 35, 3, 6, 68, -15, -28, -64, 63, 1, 11, 21, 37, -20, 8, -33, -32, 7, 58, 24, 25, -80, 8, -34, 98, -18, -33, -10, 42, 21, -44, -2, -41, 29, -9, -52, 52, -32, -74, -35, 24, -45, -35, -8, -37, 46, -24, 1, -43, -1, -13, -39, 57, -35, -72, -37, 0, -4, -22, 6, -68, -33, 0, -45, 8, 31, 26, -1, 49, -44, -54, -11, 30, -19, -11, 4, 11, -12, -47, -50, -55, -6, -12, -1),
    (-90, 9, -23, 11, 3, -40, 5, -22, 30, -35, 21, -28, -32, -47, -11, -59, -28, 12, -12, -37, 10, -23, -33, -31, 22, 10, 41, -19, -21, -23, 38, 18, 1, 32, 34, -14, 16, -38, 30, 5, 73, 37, 38, -18, -35, -30, -49, -29, -44, 70, 33, -38, -17, 22, -39, -15, 27, 22, -13, -17, -45, -2, 26, 56, -3, 5, 34, 17, -20, 26, 22, -3, 24, 41, -44, -40, -5, 15, 10, 28, 35, -10, -47, 18, 56, 12, -37, 0, 23, 39, -23, -64, -23, -6, 0, -63, 2, 25, 42, -14, -41, 41, -25, -18, -26, -16, -34, 28, -20, -28, 17, -28, 32, 65, -6, -38, 15, -18, 20, -3, -21, 35, -38, 7, -55, -22, 15, 9, 73, 4, -13, -47, 47, -66, 14, 13, -61, -6, -38, 21, -13, 0, -25, 7, -5),
    (20, -14, -33, -6, 1, -30, 36, 50, -48, 3, 15, -2, 48, -18, 46, 26, -5, -7, 40, 2, 11, -43, 36, -36, -9, -47, -27, -4, -1, 52, -9, -8, -36, 38, -17, -8, 18, 8, 24, 21, 19, -11, -2, -26, -9, 24, 49, -5, -16, 9, -3, 64, 23, -31, -35, 7, 46, 32, 54, 50, 4, 9, 38, -61, -48, -10, -8, -2, 86, -32, -41, 54, 66, 35, 6, -37, -38, 2, 5, -85, 20, -14, 5, -58, 55, 68, -74, 34, 46, 0, -37, -56, -37, -13, -1, 19, 13, -15, -42, -68, -10, 42, -41, -12, 24, 11, -81, -62, -19, -48, -51, -3, 34, -13, 6, -62, 21, 56, 17, 13, -51, -50, -27, -81, -57, -42, -13, -13, -31, -30, 47, 37, 9, -55, 22, 31, -63, -57, 39, -42, -41, -28, -13, -61, -2),
    (-21, 19, -24, 15, 19, 1, 35, -19, -14, -25, 44, 29, 1, 18, -28, 8, 6, -12, -15, 8, -22, 6, -20, 34, -11, 20, 25, -17, 10, 0, -31, 13, 14, 16, 25, -49, 13, 97, -4, 9, 8, 22, 4, -4, 14, -12, 32, -5, -60, 45, 44, -38, -11, -29, 72, -49, -6, -15, 55, -10, 11, 35, -19, 2, -21, 28, 43, -19, -25, 29, -13, -29, -14, -37, 40, -28, 9, -21, 34, -7, -10, 32, -12, -50, 12, 42, 19, -25, -42, -1, 13, 5, 57, -6, 29, -32, -9, 33, 39, -13, -33, -18, 31, 32, 23, -14, 49, -31, 28, 0, -36, 17, 5, 36, 12, 9, -39, -6, -26, -15, 46, -3, 8, -10, -3, 46, -53, -33, -46, -20, -6, -7, 7, 17, 31, -22, 7, 0, 23, 21, -46, 41, -24, -14, -5),
    (-26, 22, 27, 31, 38, 19, -5, 38, -2, 41, 49, 11, 14, 9, -13, -31, 20, -22, 12, 16, 82, -46, 24, 25, -14, 21, 44, -49, 22, -14, -68, -20, 5, -82, 16, -47, 89, 7, 7, -2, 35, 22, -44, -60, 13, -60, -15, -40, 46, -42, -56, -5, 43, 23, -55, 39, 8, 34, 17, -7, -3, -43, -48, 19, 42, -74, -1, -92, 89, 12, -63, 29, 1, -30, -54, 6, -83, -60, 35, -12, 17, -102, 10, -98, 73, 26, -39, 16, -11, -68, -14, 22, -65, 42, -17, 4, 20, -25, 5, -25, -29, 4, 14, -5, -21, -41, -41, 52, -49, -22, -2, 39, 38, -87, 21, -58, 14, 25, -20, -48, -34, -63, 15, -16, -44, 33, -25, 7, 15, -66, 46, 15, 40, 1, -20, -32, -11, -13, 51, 21, 13, 49, 15, -3, 7),
    (4, -18, 15, 54, -23, 66, -19, 28, 34, 30, -8, -36, -10, -18, 29, -52, -16, 40, -5, 4, -72, -5, 52, 32, 41, 1, 72, 19, -12, 37, -24, 33, -36, 8, -23, -6, -57, 28, 53, 22, 12, -48, 59, 7, -24, 39, 4, -21, 33, 61, 43, 19, -74, 61, -41, -28, 2, 20, 28, -66, -42, -15, -38, -16, -10, 63, 37, -5, -119, 4, -25, 4, 8, -28, 51, -52, -33, 7, 16, -3, -4, 51, 24, 21, -79, 54, -27, -37, 45, -4, 12, 4, -32, 5, -30, -9, -22, 46, -16, -12, -20, 30, 5, -29, -49, -14, 50, 47, -21, -42, -56, -23, -20, 6, 41, 0, -35, -12, 17, -61, -53, -23, -25, -21, 30, -48, -54, -24, 26, 29, 39, 13, -33, -3, -10, -17, 16, 39, -14, -44, 33, -21, -13, 3, -5),
    (13, 29, -74, 41, 12, -37, -66, 19, -53, -53, -70, 26, -36, -44, -36, 10, 2, 45, -6, -15, -59, 24, -46, 6, -33, -6, -44, -49, -17, -22, 52, -33, -23, 72, -32, -26, -56, -12, 19, -37, 10, 49, -8, 23, -27, -44, 44, -44, -15, -36, 23, 4, -48, -2, 23, -6, -69, 35, 13, 34, 43, 25, 27, 42, -47, 18, 22, 12, -1, -20, 11, 42, 10, -28, 25, 54, -28, -34, 20, 18, 46, 63, 19, 27, 10, -6, 11, 9, 0, -60, -34, -6, 45, -30, 55, 0, 71, -14, -4, -5, 1, -2, -48, 8, 6, -26, -24, -8, -27, 22, 56, 7, 0, 26, -22, 34, -9, -10, -9, 54, -38, 43, -31, 49, -76, -22, 60, -37, 39, -41, -58, -6, 14, 23, -29, 15, -7, 6, 11, 31, -21, -17, -8, 3, 8),
    (16, 18, -49, 30, 5, 63, -27, 42, 21, 71, -10, 49, 9, -2, -7, -30, 15, -9, 8, 35, 12, -1, 4, 65, 37, 55, -44, 78, 18, 17, 47, -45, 20, -28, 5, -17, 51, 38, 7, 34, -20, 54, 9, -9, 4, -6, 18, -11, 31, 39, -47, -39, -73, 78, 27, -33, 9, -22, -21, 13, -39, 27, 27, 43, 49, 26, -39, -83, -53, 100, -18, -63, -46, 15, -27, 70, -36, -27, 15, 65, 7, 12, -13, -86, 18, 11, 0, -18, 1, -42, -44, 21, 22, -16, 33, 54, -40, -5, 31, -19, -11, 38, -11, -14, 13, -25, 31, -30, -19, -15, -23, 29, -32, 45, 40, -12, -17, 12, 35, -6, 55, -30, -10, 41, -28, 19, -27, 67, -3, 55, -13, -56, -23, 45, -43, 32, -11, -40, 51, -17, 17, 5, -24, -7, -1),
    (18, 38, -26, 5, -27, 11, 15, -5, 7, 1, 70, -4, -50, 26, 30, 21, 3, 38, 47, 4, -54, -68, -42, -21, -17, -37, 46, -63, -53, -25, 18, 48, 21, -25, 17, 12, 0, -17, -4, 2, -1, -26, 34, 26, -34, -56, 38, 18, 9, 51, 23, -28, -32, -18, 54, 39, -26, -16, -6, 30, 6, -8, 54, 11, -41, 5, -2, 18, -63, -28, 23, -28, 31, 3, 66, 2, -29, -8, -7, 24, 7, -45, 1, -1, -46, 6, -4, 11, -24, -46, 45, 4, -43, 7, 16, -1, 26, 15, 54, 0, -32, -27, 23, -8, 42, -23, 28, 17, 2, -25, -3, 14, -2, 56, 53, 49, -81, 19, 53, -29, 46, -31, -19, -65, 6, 29, -36, -2, -30, 26, -4, 17, -67, 13, -15, -38, -15, -23, 8, 7, 16, -6, 23, -27, -4),
    (11, -61, -27, -15, -13, -31, -20, 3, 34, -39, 20, -10, 20, 19, -21, -35, -6, -45, 21, -15, 36, -5, 46, 27, 62, 14, 41, -39, 1, 30, 8, 15, -9, -1, -8, 4, 7, 30, -41, 48, -25, 33, 1, -10, -10, -35, 39, -21, -34, -37, 41, 41, 17, -47, 48, 10, 21, -10, -2, -1, -19, -12, -24, -22, -3, -27, -15, -21, 4, 30, 41, -19, 48, 14, -16, -22, 47, 38, 6, -16, 53, 5, -28, 15, -19, 16, -54, 27, -17, 55, -48, 22, -59, -40, 18, -4, 22, 31, 16, 36, -5, -12, 32, -47, 32, -7, 44, -40, -31, 37, -32, 41, 7, 67, -7, 55, -26, 28, -3, -6, 14, 8, -35, -18, 20, -13, 24, -10, 12, 58, 3, 18, -16, 2, -29, -21, -27, 25, -27, 45, -7, -54, 10, 19, 12),
    (21, 42, 32, 52, -41, 91, -24, -1, -1, -9, 15, 51, -4, 5, -25, -29, 37, 29, -46, -27, -12, 49, 22, 57, -45, -13, -53, 4, -55, 13, -6, 55, 55, -40, -36, -30, -6, -17, -24, 50, -65, 58, -28, 65, -6, 16, 66, 8, 37, -40, -6, 44, -10, -8, -21, 69, 13, 31, 14, 24, -11, 61, -1, -6, -17, 34, 15, 33, 61, 20, -4, 10, 38, -18, 4, 94, 4, -34, 27, 11, -31, -42, 33, -3, -15, -20, -45, -14, -36, -14, -8, -5, -40, 19, 61, 51, 64, -2, -43, 53, -42, 3, -64, -45, -1, 48, -31, 4, 43, -62, -43, -35, 61, 1, -9, 51, 43, 11, -12, 9, -8, -33, -20, -37, 55, -19, -8, -41, 22, 28, 44, -21, 34, 26, -32, 8, -42, 46, 17, -32, 37, -43, -29, 27, -3),
    (25, -45, -1, 50, -41, 40, 39, 7, -14, 29, 35, 10, -27, 44, 66, -81, 0, -116, 15, 9, -15, -47, 58, 52, 21, -32, 52, 19, -17, 27, 79, -70, 8, -87, 37, 6, 23, 6, 14, 45, -35, -41, 65, 6, -10, 12, 28, -7, 29, -111, 12, -33, 10, -56, 3, -30, 20, -39, 59, -66, -18, -6, -8, 14, -7, -13, 52, 0, -40, -28, 40, 6, -11, 23, 32, -63, -24, 13, -14, 11, -37, 3, 36, 39, -30, 26, -19, 32, -22, 14, 19, -34, 46, 16, 50, 43, -8, -10, -9, 31, 35, -1, -1, -15, -34, -32, 22, -38, 0, -4, -25, -7, -3, 36, -8, -3, -17, -14, -65, -39, -35, 7, 8, -52, -32, -10, 8, 12, 19, 24, 9, 12, -42, -25, -5, -40, 2, -44, 17, -28, 17, -71, 6, 27, -5),
    (9, -35, 39, 22, 40, -22, 45, 61, 10, -22, 58, 28, 23, 55, -46, -53, -37, -65, -52, -12, 52, -68, -33, 47, 47, -14, 38, -2, 11, -17, -5, -48, 11, -32, -11, -8, 36, -6, 13, 10, -33, 22, 14, -51, -30, -8, -21, -57, -59, -25, 14, -29, 68, -46, 19, -29, 30, -34, -9, -61, 5, 80, -12, 31, -31, -66, -48, -16, 56, -54, 0, -11, -12, 3, 20, -37, 12, -4, -2, -11, 21, -12, 48, 35, -5, 3, 10, -2, -37, 35, 4, -46, -17, -48, 35, -51, -29, -23, -58, 27, 34, -27, -6, 16, 45, 8, -30, -39, -4, -7, -24, 17, 7, 15, -38, 18, 81, -11, -8, 15, -30, -6, -49, 48, 16, -34, 16, 16, -15, -19, 39, 64, 18, 33, -37, -37, 31, -6, 17, 50, 30, -5, 35, 13, 6),
    (-16, 52, -35, -2, -12, 26, 31, 34, -5, -13, 31, 3, -19, -28, -2, 52, 15, 56, -29, 11, -5, 44, 24, -9, 21, -28, -22, -5, -10, 34, 46, 14, -37, 46, -46, -52, -36, -15, 27, -23, 2, -31, 9, -9, 1, -28, 11, -17, -33, 19, -50, 53, -48, -52, 6, 16, 18, 3, 52, 53, 14, 47, 31, -21, -52, 35, -25, -12, -49, 5, 87, 46, 10, -56, -1, 16, -21, 10, -34, 36, -4, 21, -18, -30, -36, -11, 19, 40, 40, -63, 14, 0, -38, 39, 30, 9, -7, 10, -54, 43, -12, 36, 53, 19, 18, 17, 26, 30, 7, -41, -32, 18, -28, 51, -41, 17, -44, 40, 65, -3, 28, 3, 11, 23, 2, 2, 62, -5, -24, 47, -15, 16, -13, -6, 44, -21, -25, -13, -40, 26, -8, 50, 30, -4, 6),
    (-6, -5, 8, 1, 42, 4, 14, 43, -12, 6, -4, 24, 33, 15, 40, -17, -16, 28, 15, 48, 18, 50, -53, -18, -9, -86, 38, 14, 37, -7, 53, -12, 18, 32, -61, -59, 26, -54, -55, -5, 1, -62, -41, -13, 11, -9, 53, 2, 40, 1, -52, 59, -16, 48, -33, 10, 7, 14, -46, -8, -43, -23, 11, 53, 9, -13, 25, 37, -9, -19, -43, -37, -23, 38, 22, -44, 12, 18, 29, -55, -20, -49, -47, 19, -11, -21, -19, -31, -16, -9, -61, -7, 5, -5, -26, 9, -34, 25, -34, 32, -53, -8, 50, 22, -5, -74, 19, 31, -21, 3, -33, -6, -1, 36, -52, 7, 22, 12, -23, -18, -61, 1, -15, 33, -72, 14, 28, 8, -40, 42, -65, 6, -16, 25, 39, -35, -37, -39, 24, -6, -32, -65, -24, -6, 0),
    (-84, 21, -31, -32, -72, 58, -43, -10, -52, -49, -8, -27, 3, -49, 11, 47, -15, -28, 18, -8, -13, -61, 6, 0, -1, -14, 52, -19, 36, 18, -14, 2, 26, 40, -15, 21, -3, -28, -21, 23, -27, -7, 37, 20, -1, 9, -33, 4, -37, 62, -14, -14, -53, -11, -31, -11, -58, 5, -68, 59, 35, -20, -28, 34, -54, 60, 0, 38, -91, 19, -45, -33, 51, 18, -23, -69, -21, -53, 50, -11, 28, -9, 1, 16, -51, 5, 7, 57, 8, -13, 37, 49, 3, 48, 25, -15, 0, 39, -8, -13, -20, -4, -3, -4, -6, -39, 2, 18, -30, -4, -30, 2, 43, 66, -41, 1, -59, -1, -22, 11, -41, 78, 20, 8, -52, -47, -3, -4, 16, 34, -5, -5, -45, -11, -28, -60, 30, 28, 48, 13, -13, -37, 19, 31, -3),
    (-29, 44, 11, -9, -78, 0, -10, -11, -16, 32, -44, 30, 9, -23, 4, 1, -4, 40, -3, 13, -33, -21, -37, 13, -49, 32, 30, 94, 16, 25, 33, -4, 28, 4, 19, 12, 5, 5, -9, -8, 17, 37, -33, 17, -25, -22, 49, -34, -27, 8, -22, 19, 5, 37, -25, -20, 24, -18, -60, 25, 7, -37, -17, -5, 30, 3, -10, 14, 14, 27, 4, -32, -32, 61, 2, 53, 41, -46, 18, 30, 78, 21, 2, 15, 13, -44, -3, -11, -46, 64, 1, 31, -35, -28, 14, 21, -16, -17, -50, 23, 12, 6, -70, -16, -34, -19, -4, -8, 30, -56, 17, -5, 29, -8, -17, 47, 44, 14, 24, 37, 16, 33, 19, -39, -31, -59, -28, 32, 65, -27, 0, 26, 30, 5, 7, -46, 19, 28, 21, 6, -27, 0, 56, -44, -2),
    (29, -23, 13, 26, 67, -4, -17, -22, 22, 40, 53, 12, 0, -49, -10, -83, 40, 17, 34, 49, 28, -9, 29, -36, -47, 85, -1, -1, 13, 21, 13, -49, 23, 38, 39, 48, -13, -12, 36, 28, -54, 46, 22, -37, 12, 30, -19, -17, 65, -42, 12, 68, 1, -62, -13, -4, 33, 38, -1, 21, -50, 8, 73, -10, 102, -31, 9, 36, -39, -10, 56, -3, -39, 95, -15, 57, -6, 31, -6, -25, 5, 1, 20, 9, 0, 40, 12, 7, -60, 51, 14, -23, 4, 32, 12, -1, 7, 14, -36, 47, -27, 1, 35, 56, -45, 34, 3, 7, -36, -23, 50, 33, 69, -7, -37, 29, -20, 5, -25, 21, -29, 50, 23, 35, -27, -22, 63, 25, -2, -32, -18, -45, -8, -35, 16, -35, 12, 1, -38, 8, -14, 39, -47, 28, -6),
    (18, -43, 8, -16, 50, -22, -17, -36, -5, 48, 20, -6, 43, -1, -22, -59, 61, -31, 25, -29, 63, -31, 20, 45, -20, 26, -36, -8, -27, 18, 32, -57, 47, -7, -28, -14, -33, -17, 7, 5, -9, 50, -17, -8, -33, 30, 0, -16, 31, -34, -2, 25, 11, -68, 2, -42, -4, -9, 38, -2, 30, 33, 6, 7, 52, -33, 84, -12, 45, -89, -25, 25, 0, -19, 65, -42, -23, -10, 22, -39, 55, -35, 58, -51, 4, -50, -36, 8, -15, -32, 61, -36, -22, -48, 32, -93, -12, -7, -21, 16, 19, -45, 47, -36, 0, -15, 15, -35, -20, 43, -10, -12, -40, -10, 58, -27, 39, -4, -9, 6, 43, -24, -25, 31, -36, 47, 17, -38, -11, -5, 43, -8, -23, 9, -27, -18, -23, -10, 17, -6, 46, 17, 43, -51, -4),
    (18, 15, 28, 37, 58, -47, 56, 54, 35, 38, 38, 20, 44, 7, 58, -33, 2, -5, 24, 40, -16, 5, -23, 29, 5, 35, 12, 50, 78, 37, -19, -11, -25, 19, 2, -5, -31, 54, 21, -11, -39, -44, -45, -38, 50, -23, -14, 11, 15, 23, -58, 69, 32, 7, -38, 53, 7, 39, 12, 59, 60, -36, 52, -38, 0, 69, -8, 45, -31, 103, -52, 39, 15, 61, -2, 58, 26, -2, 57, -52, -33, 38, 14, 34, -49, 10, -8, 39, 30, -13, -8, 38, 19, -42, -4, 42, 25, -22, -10, 38, 4, -16, -18, 27, -44, 14, 20, 23, -30, -32, 27, 21, 40, 52, -75, -24, -14, 20, 33, -61, -37, 29, -55, -2, -90, -51, 29, -12, -22, -5, -54, -11, -43, 7, -34, 38, -26, 3, -91, -33, -46, -17, 50, 34, 7),
    (27, -19, -20, -40, -44, -69, 7, 31, 31, 7, 16, 9, -60, -13, -8, -8, 37, -46, -43, 21, -38, -15, 77, 41, 5, 21, -38, 23, 13, -29, 10, -20, 48, -32, 33, 51, -37, 8, -17, 12, 22, 0, -33, 21, -12, 37, 0, -31, 2, -10, -6, 19, -25, -2, 77, 11, -40, 35, -17, 41, -73, 44, 14, -61, 62, -13, -53, 49, -25, 69, 56, 6, 28, 79, 16, 20, -46, -17, 33, -37, -3, -29, -33, 19, -30, 29, 62, 57, 15, 60, -20, 70, -77, 29, -4, -13, 5, 37, 35, 22, 11, 20, 28, -32, 20, 8, -9, 31, -56, -22, 22, -39, 30, 31, -4, 15, -46, 24, 6, 23, 39, 45, 20, 38, -51, -13, 16, -15, 34, 48, -23, -30, -24, 25, 11, -32, 41, 42, -10, 34, -30, -50, 33, -48, -3),
    (-30, -17, 35, 14, -25, 39, 5, 9, -4, 13, 12, -36, -42, -14, 5, -5, -21, 7, 16, 24, -23, -34, -13, 36, 40, -10, 67, 3, -45, 12, 20, -41, 20, -62, 32, 30, -20, -18, 28, 12, -25, -10, -33, 18, -17, 7, 26, -50, -19, -15, 27, 54, -8, 1, 22, 4, 30, 48, 32, -30, -23, -28, -30, -35, -36, -17, 52, -31, 11, 38, 26, -48, 28, 0, 98, 3, -45, 25, -7, -76, -23, -27, -19, -16, 10, 68, -10, -23, -46, 18, 60, 33, -50, 23, 15, -86, -22, -36, -23, 11, 26, 8, -83, -17, 17, 16, 31, -11, -3, 4, -16, 10, -7, -16, 57, 24, -5, -6, -16, 25, 5, 43, 52, -2, -23, -42, -32, -52, 3, -5, 2, -15, -14, 12, 40, 13, -36, 52, -16, -14, -46, 36, -16, -55, -5),
    (-28, -18, -39, 17, -44, 22, -57, 12, -16, -27, -36, 29, 42, 1, 58, -59, 6, 4, -4, 35, 13, -36, 3, 8, 31, -14, 38, -52, -26, -12, 18, -2, -1, 12, -11, 4, 45, 27, 31, -53, -16, -8, 57, 18, -6, 34, -53, -41, 67, 23, -18, -16, -3, 36, -37, 61, -23, 70, 0, 42, -7, -62, -6, -6, 20, 45, -30, 20, -13, -45, -52, 42, -7, 67, -28, 69, -27, -38, 48, -30, 35, -2, -27, -30, -22, -7, -5, -18, -36, 29, -29, -16, 12, -28, 24, -7, 2, 10, -19, 33, -64, -18, -1, 25, 28, 5, 32, 67, -51, 57, -24, 29, 17, 19, 1, 13, -77, -16, 35, 50, -28, -3, -14, 63, -37, 27, 4, -10, 26, -6, 36, 39, -38, -51, 51, 64, 13, 3, -29, 57, 12, 1, 24, 15, -3)
  );
  ----------------
  CONSTANT Layer_4_Columns    : NATURAL := 16;
  CONSTANT Layer_4_Rows       : NATURAL := 16;
  CONSTANT Layer_4_Strides    : NATURAL := 1;
  CONSTANT Layer_4_Activation : Activation_T := relu;
  CONSTANT Layer_4_Padding    : Padding_T := same;
  CONSTANT Layer_4_Values     : NATURAL := 24;
  CONSTANT Layer_4_Filter_X   : NATURAL := 3;
  CONSTANT Layer_4_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_4_Filters    : NATURAL := 24;
  CONSTANT Layer_4_Inputs     : NATURAL := 217;
  CONSTANT Layer_4_Out_Offset : INTEGER := 3;
  CONSTANT Layer_4_Offset     : INTEGER := -1;
  CONSTANT Layer_4 : CNN_Weights_T(0 to Layer_4_Filters-1, 0 to Layer_4_Inputs-1) :=
  (
    (-7, 24, -9, -19, -10, 6, 0, 9, 13, 30, 11, -15, -11, 5, 35, -20, -23, -54, -5, -2, -14, -22, 22, -46, -30, 47, 40, -10, 42, 17, 18, 50, 24, 37, -22, 15, 31, 34, 29, 17, -44, -42, 27, 27, 29, -13, -26, -5, -21, 33, 45, 44, 4, 19, -10, -11, -3, 38, 18, -8, 6, 16, 62, -13, 3, -7, 19, -12, -9, -13, 43, -3, -35, -39, -20, 12, -21, -30, 27, 29, 7, -50, -22, 5, 7, 2, -63, -19, 13, -11, -25, -15, 11, -50, 1, 4, -46, -14, -8, 27, -20, 17, 30, -14, 25, 2, -34, 21, -38, 10, -41, -23, -26, 54, 22, -21, -21, 30, 4, -42, -56, 5, 15, 14, 31, 64, 11, -1, 7, 9, -25, 24, 31, 29, 19, -54, -42, 30, 15, -3, -13, 32, 43, 22, 34, 20, 34, 9, 7, 19, -23, -34, -16, -37, 1, 4, 3, -37, 19, -32, 41, 33, -30, -38, 28, -4, 5, 24, 3, -74, 20, 64, -33, 37, -32, -11, -5, 19, -51, -22, 11, 21, -17, 7, 15, -14, 21, 10, -20, 9, -47, -10, -39, -77, 24, 12, -2, 27, -26, 11, -20, -49, 2, 0, -25, -4, -73, 33, -24, -20, 27, 43, -23, 24, -32, 17, -4),
    (-9, 42, 2, 2, 10, 35, -43, -12, 36, -11, 7, 27, 27, 19, 56, -17, 12, 19, 25, 46, 54, -1, 25, 59, -18, -24, 3, 5, -33, 8, -64, 45, 15, 7, -21, -31, 14, 1, -21, -46, -11, 41, 32, -10, -25, -25, 7, 32, -28, -68, -58, -3, -3, -4, -37, 30, -67, -27, 5, -21, -5, -9, 2, 21, 24, 12, 1, 13, 13, -35, -18, -9, -9, 26, 24, 4, 6, -16, -15, 19, 13, 12, 15, 20, 7, 28, 30, 18, -4, -47, 24, 16, 31, 57, -3, -30, -43, 17, -33, 8, 40, -23, -18, -2, 15, -22, -23, -31, 15, 31, 21, -11, -11, 7, -1, -9, 36, 20, -29, -13, -59, 18, -2, 31, -28, 22, 8, 5, -8, 13, -25, 5, 38, -5, -40, 4, -32, 34, 2, 9, 16, -3, -31, -15, 50, -9, 13, 0, 11, -2, 19, -38, -38, 21, -11, -64, -47, 10, -42, -4, 22, -21, -52, -18, -2, -30, -45, -19, -6, 20, 28, -22, -28, -30, 9, -10, 15, -33, 24, -28, -12, 5, 12, -15, 2, -15, -19, 23, 29, -18, -34, -10, 9, -21, -9, 36, -31, -25, 31, 6, 19, -37, 5, 18, 32, 2, -36, 14, 7, -64, -39, 10, 13, -41, 17, -25, -2),
    (-52, 8, 59, -11, -61, -18, 10, 38, -54, -16, -46, -38, -4, -52, -50, 32, -77, 6, 0, -32, -6, 4, -11, 28, 16, 43, 63, 31, -32, 11, -33, 8, 15, 8, 4, -63, 2, -50, -31, -9, -32, 0, 10, 11, 17, 7, -36, 19, 10, -10, 6, -21, 18, 37, -6, -23, -12, -51, -24, -66, -34, 5, -46, -45, 1, -49, -32, 21, -2, -37, 21, -25, -50, 21, 6, 34, -4, 11, 3, -46, -20, 24, 8, 35, 49, 38, -6, -18, -40, -37, -11, -19, 37, 32, 16, -2, 15, 16, 42, 4, 16, -11, 43, 3, 28, -12, 43, 15, 21, -24, 39, -23, 21, -9, 6, -22, 11, 22, 25, 52, 53, -30, -61, 3, 1, -52, -7, 32, -4, -19, 5, 9, 19, -9, 22, 8, 39, -38, -33, -7, -31, -39, 33, 4, 8, 13, 59, 13, 10, 28, 33, -9, 34, 2, -30, 11, 44, 17, -65, -69, -15, 12, -2, 26, -18, 4, -10, -7, 53, 6, 24, 13, 34, -41, 12, 1, 43, -27, -34, 50, 30, -34, -28, -42, 44, 62, -16, 23, -59, -34, 28, 15, 36, -8, -19, 12, 11, -15, 45, 24, -30, 26, 11, 24, 16, -17, -31, -26, 13, 51, 12, 13, -63, -48, -2, -24, -6),
    (6, -6, -9, -9, -8, 5, 1, 2, -78, -26, 15, -25, -20, 44, -21, -30, -1, -59, -12, 61, -34, -6, 24, -51, -49, -13, 26, -15, 6, 17, -24, -9, -35, -21, 7, -42, 26, 67, -6, 48, 44, -43, -15, 35, 30, -13, -34, -36, 64, 26, 29, 11, 23, 32, -23, -27, 9, -32, -23, -5, -11, 0, -61, -12, 52, -7, 58, 9, -7, 1, -36, 11, -11, -36, -15, -26, -2, 14, 41, -4, -33, 23, 52, 27, -10, 8, 9, -14, 10, 19, -30, -7, 59, 22, -7, -28, -49, -33, 10, 24, -43, 9, -70, 35, 27, 3, -21, 11, -37, -23, -7, 15, 12, -2, 19, -12, 27, 16, 6, -8, 40, 0, -30, -9, -10, -36, 37, -8, -2, -48, -27, -6, -39, -42, -18, 41, 3, -14, 5, -54, -10, -9, -7, -36, -37, 66, 12, -17, 16, -35, 8, 28, 2, -9, -5, 80, 24, -47, 1, -19, -51, 0, 11, -7, 45, 14, 14, 44, -62, 6, -19, 62, -26, 26, -4, 44, -16, -53, -18, 41, -28, -31, 11, -19, -35, -32, 42, -22, 30, 37, -29, 35, 35, -30, -1, 48, -32, -33, 30, 6, -73, 6, -45, -63, -6, -6, -22, 25, -21, -4, -59, -6, -29, -14, -17, -40, 12),
    (2, -17, -12, 56, 34, 22, 11, 25, 23, -37, 23, 62, 11, 4, -11, 10, 39, 69, 52, -31, 21, -2, -28, -1, 31, 1, -19, 8, -9, -1, -16, 13, 49, -16, -34, 39, 21, -12, 20, 41, -10, 49, -26, -26, -6, -29, -35, 47, -12, -37, -36, 0, 9, -39, -15, -3, -11, -14, 13, -31, -44, -6, -47, -12, -31, -25, -67, 3, -6, -15, -16, -7, -17, 59, 23, 29, 20, 19, 45, -27, 100, 19, 26, 62, -2, -23, 22, 13, -16, 67, 48, 21, -8, 8, -21, 27, -25, 46, 4, 26, 21, 38, -23, 23, 76, 28, 22, -53, -7, 8, -3, -18, 37, 8, -35, 31, -37, -47, -42, 5, -52, -16, -9, -56, -15, 19, -8, -22, 6, -36, 9, -59, -41, -42, -19, -51, -8, 35, -32, 37, -4, -39, -28, 0, -69, 2, 26, 21, 0, 19, -12, -67, 61, -47, 12, 16, -12, 7, -30, 39, -8, -42, -37, -21, -32, 28, -45, 11, -62, -3, 16, -12, -22, 20, -1, -17, -14, -28, -27, -54, -8, 57, -22, 31, -39, -19, -50, -11, -38, -26, 9, -66, 13, 11, 13, 10, 29, -76, 8, -5, -33, -4, -27, -9, -26, 48, 6, -57, 49, -12, 4, -14, -16, -15, 7, -50, 7),
    (39, 21, -2, 0, -26, 41, 18, -21, -26, -1, 6, 36, 23, 2, 28, -21, 6, 54, 18, 8, -8, 0, 34, 7, 30, 9, 29, -6, -5, -30, 29, -3, 43, 15, -34, 13, 41, 12, 6, -7, 20, 6, 4, -7, -6, 35, -13, -4, 28, 24, -22, -28, -7, -73, 3, -41, 32, -8, -10, -1, 9, -18, 3, 42, 18, 31, 16, 3, -13, 21, -7, -19, -7, -41, -14, 25, 2, 55, -44, 18, -49, 37, 16, 5, 13, -8, 11, -24, -26, 25, 54, 13, 37, 9, 38, 11, -15, -45, -27, 23, 7, 17, 21, -13, -29, 43, 32, -15, -36, 30, -36, 23, -52, 23, -35, -16, -51, -55, 8, -2, -1, -10, 20, -2, 5, -45, 25, -32, -65, 12, -17, -23, 3, 55, 23, -12, 1, -35, 1, -12, -32, -5, 9, -29, -101, -34, -33, 64, 10, 9, -24, 6, -15, 44, -5, 17, 16, 20, -11, -11, -49, -43, 48, 50, -5, 7, -22, -29, -33, -42, -30, 22, 31, 35, -12, -41, -28, -8, 11, -27, 23, 14, -22, -21, -46, -31, -10, 26, 19, 14, 27, -45, -28, -22, 20, -5, -33, -13, -10, -46, -57, 17, 6, 1, 21, 36, -1, -16, 36, 24, -14, 8, 20, -26, 35, 12, -2),
    (1, 51, -16, -36, -26, 23, 15, -19, 18, -20, 41, 91, -4, -1, -32, 61, -54, 33, -22, 36, 53, -5, 21, -6, -25, -11, 21, 59, -56, -18, 10, -58, 41, -5, -18, 46, -24, 27, -20, 37, -23, 16, 9, 31, -21, -32, -25, -11, -21, -2, -20, 4, 36, -8, -31, -27, 52, -34, 25, 29, 17, -19, -6, -30, -11, 19, 28, -1, -52, -20, -42, 6, 19, -19, 4, -2, -12, -40, 8, 27, -63, 30, -21, 1, -41, -26, 28, -30, -24, -14, -10, -10, 19, -58, 6, 30, 34, -33, -22, 15, -58, -81, -11, 0, 42, -46, 5, -21, -35, 24, -38, 0, 83, 31, -4, -50, -1, -13, 0, -28, 45, 10, 7, 57, -14, -67, 26, 30, -13, -10, -53, 14, -1, -12, 16, 24, 15, 11, 46, -31, -12, 24, -33, 17, -8, -4, -8, 4, 9, 37, 8, 27, 26, -15, -21, -5, 12, -16, -4, 17, -29, -22, 0, -14, 56, -10, 6, 16, 8, 26, 17, 25, -33, -33, -14, -30, -16, -41, -53, 50, -13, 21, 40, 27, 18, 24, -20, -28, -7, 1, 14, 9, -14, 5, -30, 63, 33, 40, -26, -16, -16, -3, -51, 17, -26, -3, 17, 3, 9, 29, 54, 9, -22, 35, 15, 60, -3),
    (-8, 37, 8, -4, 20, 25, 35, 17, 20, -28, 23, 21, 34, 54, 13, 4, -3, -12, 13, 35, -12, 34, 41, -38, -20, 1, 37, -19, -2, 17, 1, 60, 13, 22, 32, 29, 27, 13, 34, 28, -16, 33, 40, 17, 18, 32, 20, 7, -24, 34, 28, -5, -20, 18, 6, -26, -1, 26, 5, 38, 54, 40, 5, -22, -67, -17, -2, -3, 25, 7, -35, -33, 32, -34, 1, -31, -18, -17, 9, 23, -32, -20, 23, 30, 18, 15, 9, 17, 4, -28, -60, -12, 6, -18, -16, -64, 78, -28, 33, -55, -21, -22, 29, 0, -32, -8, -4, 4, 27, -10, 25, 35, 36, -26, -42, -2, -29, -53, -35, -37, -34, -11, -52, -26, -23, -41, -28, 10, 4, 11, 15, 13, -51, -17, -20, 46, -12, -73, -6, -35, -4, -40, -36, -18, 35, -36, 9, -10, -21, -32, 29, -40, -46, -42, 31, 9, -47, -16, 17, 39, 42, 69, -29, 2, -29, -29, 8, 0, 67, 43, -8, -54, -4, -71, 10, 53, 35, -34, 10, -3, 23, -39, 37, 27, 45, 7, -16, 2, -24, -31, -14, -17, 46, -32, 10, -4, 7, -20, -24, 22, -9, 19, -16, 58, 15, -39, 5, 41, 33, -25, -58, -29, 22, -18, 6, -16, 9),
    (9, 68, -24, -37, 36, 3, -30, -4, 21, 8, 35, 16, -4, -37, 38, 36, 32, 18, 16, 28, -51, 14, -44, 32, -71, 56, -7, -50, 14, -21, -22, 51, 28, 0, -5, -1, 4, -36, 33, -14, -16, 13, -37, 18, -35, -32, -30, 11, 5, 27, -41, -11, -36, -25, -13, 1, -6, -46, -24, -42, -50, 12, 13, 17, -48, -9, -37, 11, -12, -25, 23, 16, 53, -10, -30, -19, 31, -22, -12, 0, 11, 20, -18, -3, 27, -16, 81, 15, 59, 14, -55, -33, -38, -22, 28, -6, -31, 42, -24, -40, -5, -12, -48, 22, 31, -24, -54, -42, -45, 15, -16, 29, 21, -7, -41, -22, -12, 14, -35, 11, -22, -7, 14, -12, -33, -24, -59, 33, -16, -6, 19, 9, 9, -31, -26, -34, -14, -18, 32, -39, 6, 9, -11, -29, 16, 14, 17, -56, -1, -16, 1, 32, -21, 43, -7, -20, -12, 1, 56, 20, 35, 4, -23, -20, 43, -18, 16, 42, 31, 54, 49, -17, -10, 24, -20, 17, 33, 33, 7, -20, 32, -8, 16, -13, 29, 11, 34, -16, 19, 4, -16, 12, 8, -15, -12, 40, 1, 26, -19, 7, 9, 8, 25, 58, 5, -23, -29, -15, -35, 1, -27, -21, -8, 2, -3, 19, 2),
    (12, 15, 29, 75, -12, 9, -27, -18, -22, -47, -16, -37, 14, -35, -42, -3, -42, -60, 20, 37, -4, -12, 21, -36, 24, -38, 29, 28, -5, 4, 1, -23, 2, -1, 4, 42, -30, -37, -48, 37, -5, -9, 12, 2, -59, -3, -12, -13, -23, 22, -10, -36, 3, -37, 44, -38, 19, 23, 10, 11, -19, -43, 1, 7, 103, -17, -41, -41, -8, -11, -33, -14, 13, -16, 7, 44, 11, 33, -4, 41, 1, 1, -23, 17, 7, 18, 16, -22, 27, -25, 47, 14, 17, 73, 42, 51, -2, -10, -2, -8, -2, -2, 17, 40, 2, 22, -1, 21, -16, -10, 55, 16, 61, 39, 62, 11, 41, 27, 20, 59, -13, -45, -81, -75, 10, -48, -13, 0, -53, 46, 2, -29, -9, -28, 60, 2, -41, -54, 6, 1, 12, -32, -49, 5, 8, -30, 9, 1, 15, -2, -24, 19, -3, -22, 7, -17, 12, -34, -29, 20, 26, -41, 12, 30, 27, -5, 28, 33, 21, -6, 23, 10, -21, 3, 32, 58, 8, 9, -4, 9, 48, -20, -13, -33, -34, 26, 39, -8, -33, 6, -29, 36, 7, -17, -8, -40, 22, -57, -4, 28, -24, -4, -21, -24, 13, -9, -18, -35, -23, -20, -12, -2, -33, -12, -26, -59, -7),
    (20, 22, 56, 15, -69, -27, -23, 10, -35, -4, -46, -9, -44, -2, -53, -21, 8, -1, -13, -42, -16, -52, -57, -48, 28, 42, -4, 49, 20, 19, 8, 27, 3, -40, -19, -18, -34, -16, -52, 5, -14, -17, -13, -49, -27, 0, -37, 15, 2, -7, 64, -3, -26, 53, -43, -51, 56, -5, -19, -30, 24, -28, 14, -67, 30, -7, -46, -43, 15, -47, 30, 10, -105, 54, -5, -19, -43, -15, -20, 72, 1, 17, -40, -46, 22, 0, 37, 10, -69, 4, 1, -17, 4, 32, 16, 22, -22, 9, 12, 8, 25, 16, -47, 11, 13, -12, 17, 8, -19, 8, 41, 3, -75, -2, -35, -56, 37, 25, 28, 34, -17, 62, 81, -25, 38, 44, -16, -6, 31, -17, -10, 29, -18, 5, 61, -21, -20, 20, -20, 23, 44, -10, -29, 28, -35, -43, -51, 21, 19, -7, -29, -23, -41, 27, 19, -6, 54, -33, -7, -46, -26, -17, 20, -15, 6, 12, -23, -21, 5, -48, 30, 11, 22, -17, 38, 0, 43, -4, 30, 3, 30, -38, -16, -31, 26, -36, 23, -28, 19, 13, 37, -53, 13, 49, 54, 18, -12, 40, 37, -9, 6, -15, 3, 43, 2, -9, -1, -7, -16, -21, -22, 26, -21, 39, 6, -16, -2),
    (-33, 17, 27, -28, 12, 8, 29, -82, 32, 45, 23, -41, 42, 40, 15, -6, -65, -82, 8, 29, 22, 13, 1, -37, 23, -17, 3, -36, 8, -60, 37, 8, -30, 63, -15, -10, 46, -11, -7, 64, 13, -39, 33, 34, 3, 32, 22, -16, -14, 34, 28, -64, 40, -51, 49, -33, -36, 53, -28, -33, -9, -29, -19, 27, 29, -7, -14, 17, 8, 25, 30, 9, -6, -18, -10, -27, 9, -37, -17, 29, 14, 3, -31, 14, -6, -17, -19, -6, -8, -12, 15, -9, -22, 8, -10, -24, 23, 12, -46, -19, 22, -52, 48, 9, -20, 26, 6, -31, -14, -19, -28, 2, 0, 10, 30, -17, -29, -34, 11, 18, 43, 0, -13, -15, 38, -47, 54, -3, 16, -16, -38, 10, 12, 5, 0, 9, 29, 41, 41, -5, -28, 12, 34, -11, -17, -5, -7, -2, 35, -21, 10, -3, -29, -25, -24, 27, -20, -1, 1, -22, -51, -9, -18, 30, 2, -17, -34, 27, -1, -33, 4, 29, -36, 15, -1, 29, -31, 11, -11, 26, 6, 20, -29, -24, -7, 4, 24, -9, -9, -12, 4, 42, -3, 11, -47, 39, -12, -20, -28, 5, -75, -1, 32, -22, -6, -18, -23, 9, -33, -7, 25, -18, -2, 6, 31, 0, -9),
    (-32, -31, -15, -50, 19, 2, -56, -20, -4, 12, -35, -42, -25, 20, 25, 6, 63, -23, -12, 17, 6, -42, -48, -24, 3, 8, -8, 5, -28, 1, 6, -2, -21, -40, -20, -15, -4, -25, -33, -19, -24, 16, 40, 32, -21, 9, 31, -66, -1, -32, -7, -47, 9, -33, 59, -20, -86, 11, -16, -37, 56, -28, -14, 0, 9, -6, 13, -12, 3, -16, -28, 3, 3, -13, 7, -16, 48, -11, -15, 35, 21, 16, 31, -20, -30, 17, 68, 49, 7, -10, -26, -19, -39, 32, 6, 20, 13, -20, 31, 27, -46, 23, 23, -7, 32, -50, -13, -38, 17, 35, -10, 56, -2, -34, -7, -50, -44, 13, 17, -3, 1, 2, 50, -10, 11, -21, 24, 10, 41, -25, 36, -25, 16, -22, -46, -35, 7, -42, 2, -21, -22, 19, -28, -47, -17, -36, -13, -22, 30, -33, 60, -30, -41, 22, -35, -19, 44, -28, -50, 4, 25, 7, -7, -30, -4, 10, -12, -4, -17, -5, -37, -21, 12, -9, -2, 36, 10, -2, -45, 23, 20, -48, -13, 11, -29, -19, -9, -56, 27, 34, 26, -39, 34, -11, -4, -7, 22, -5, 9, 16, 17, -15, 18, 18, -3, -37, 23, 0, 4, -6, -59, -58, -6, -15, -33, 1, 0),
    (-35, -16, -40, 9, 19, 11, 0, 21, -54, 17, -15, -15, 9, 14, -17, 24, -24, -45, -25, 37, 62, 21, -25, 13, 10, 18, 19, 9, 11, 36, -19, 46, -10, 5, -16, -19, 7, 43, 8, 16, 36, -65, 48, 18, 32, -20, 2, 3, -46, 4, 31, 9, 3, -3, -28, 5, -10, -30, -15, 11, -24, 37, -5, 57, 19, -67, -15, -32, 18, 22, 13, 4, -28, 11, 4, 4, 18, -8, 14, 38, -24, -24, 10, -11, 2, 36, -6, 46, -2, -38, 27, -16, 39, 16, -27, -10, 7, 13, 39, 28, 4, 17, -47, 25, 40, -42, -26, 30, -21, 0, 30, 20, -15, -1, 39, 11, 32, 66, -45, 69, -7, 41, -28, -27, -30, -9, -55, 41, 21, 23, 20, 12, -13, -28, 18, 5, -34, 16, 2, -29, -14, -16, -29, 22, 0, -43, 23, -8, 22, 16, 34, 5, 28, 36, 46, 15, 38, -12, 13, 23, 18, -8, 29, 38, 8, 10, 29, 4, 50, 39, -31, 36, -14, 0, 11, 38, 5, -9, -24, -23, -12, -56, 1, 80, -17, 14, 52, -3, 16, 39, -50, -11, -16, -18, 0, -67, -55, -50, -39, 22, 17, 17, -15, -18, -24, -77, 32, 23, -38, 38, -12, -54, -8, -23, -14, 29, 4),
    (-69, -11, -15, -6, 43, 48, 11, -44, -41, 5, 19, 27, 44, 25, 3, 12, -66, -3, -23, 47, -17, 10, 53, -36, -45, 41, -30, -35, 41, 25, 8, -6, 4, 16, 23, 18, 2, 6, -10, 77, -29, -31, 33, 34, 21, 15, 43, -33, 35, 59, 4, -8, -25, 4, 26, 23, 5, 29, -61, 31, -4, -16, -11, 51, -35, -21, -37, -8, -19, -15, -52, -25, -47, -32, 10, -8, 33, -19, 15, -62, -34, 15, 6, -10, 56, -6, 1, -24, -31, -9, -22, 20, -18, 5, 26, -49, 53, -12, 44, -32, -18, 0, 30, -4, -7, -2, 28, -15, -10, -1, -20, 22, 27, 46, 47, -8, 24, 9, 9, 25, 71, -5, 3, -3, 21, 0, 44, 3, 16, 30, -3, 5, -3, -47, 17, 16, 43, 41, 35, -46, -3, -7, -2, 1, 0, -40, -47, 27, 11, 13, 6, 14, -49, -25, 21, 0, 7, -24, -11, -36, -4, -3, 25, 37, -36, 30, -2, -8, -26, -17, -25, 5, 33, 13, -32, 2, 21, -3, -19, -14, 33, -30, -16, -34, -32, 9, 32, 22, -12, -9, 44, 23, 4, -32, 8, 3, -52, 23, -8, -7, 28, -33, -24, -1, -4, -19, -30, -4, -70, 49, -33, 2, -17, 12, 2, 20, -8),
    (-46, -53, -35, -25, 30, -67, -30, 20, -2, 24, 13, -42, -25, -4, 51, 48, -54, -53, -39, 32, 16, 36, -29, 15, -9, -6, 25, 29, -36, 2, -17, 51, 16, -22, -30, 20, 12, 16, 38, -35, -20, 38, -16, -7, 33, 22, 4, -18, 40, 29, 46, 53, -36, -1, -14, -51, -1, 10, -15, 13, -20, 28, 35, -46, 41, -8, -5, -28, 15, 22, 35, 30, 26, -21, -31, 17, 25, -21, 0, -40, 10, -18, 45, -19, 7, -16, 34, 0, -15, 14, -6, -11, 1, 16, -42, -11, 26, -21, -34, 10, -8, 28, -26, 27, 60, 13, 34, -17, -45, -29, -35, -34, 77, -31, -41, -4, 9, -29, -12, 9, -8, -21, 0, 14, 12, 19, 5, -39, 50, -28, 16, -31, 12, -5, -13, -34, 25, -3, 21, -43, 26, -9, -4, 5, 28, -9, -30, 18, 0, -2, -8, -7, 10, 15, 25, 5, 38, -7, 40, -12, 69, -29, -42, 19, -20, -26, 23, -4, 43, -66, -38, -22, 38, -28, -55, -13, 22, 20, -12, -1, -6, -18, 0, -41, 1, 9, -22, 19, 5, -54, -33, -4, 25, -64, -15, -31, 34, -38, 27, 5, 14, 38, -2, -27, -22, -13, 9, -35, -5, -27, -46, -32, -29, -47, 36, 37, 5),
    (26, -35, 23, 15, 45, 5, -53, -30, -10, 8, -17, -47, -1, -16, -10, -2, -2, -30, 8, 48, -22, -15, -31, -27, -23, 29, 43, 16, 32, 20, -12, -64, -24, 36, -29, -15, -3, -29, -40, -12, -22, -24, 19, 6, -9, -57, 42, -45, 27, -25, -36, 14, -37, 52, 15, -54, -57, -26, -10, 34, -1, -30, -36, -22, -36, -35, -16, 4, -36, -27, -23, -10, 11, -4, 37, -32, 32, -10, 27, 0, 20, 36, -25, -19, 44, -1, 23, 36, -6, -17, -4, -35, 38, 5, 13, -6, -38, 8, 34, -38, -23, 2, -21, -44, -42, 35, 17, 32, -1, 1, 6, -22, 17, 14, 57, -2, -34, 37, 14, 0, -56, 22, -8, -3, 48, 9, -48, 3, -80, -20, -11, 28, -6, -11, -30, -36, -73, 15, 35, 70, 52, -35, -17, 9, -23, 13, 15, -30, -42, 16, 29, -36, -43, -34, -14, -1, 33, 9, 21, -9, -65, 18, 4, 3, -11, 28, -10, -34, 1, 51, -28, -29, 29, -18, 33, 4, 17, -1, -33, -37, 50, 19, 52, 1, -20, 23, -19, -27, -1, 32, 32, -18, -20, -9, -9, -38, 28, 15, -11, 10, 35, 47, -30, -12, 38, -12, -9, 9, -23, 41, 32, -8, -3, -19, -10, -32, -5),
    (1, -19, 33, 27, -8, -45, -41, 64, 14, -29, -31, 45, 5, -33, -45, 29, 32, 68, -22, 9, -11, -23, -18, 47, 39, -14, 19, 21, -31, 16, -45, 14, 34, -34, 16, 57, -27, -18, 10, -40, -46, 23, -5, -21, 8, -47, -40, 28, -40, -60, -39, -8, 27, 35, -24, -14, -31, -24, -5, 32, 35, 33, 36, -34, -16, 25, -19, -38, -58, 2, 17, -30, -56, -66, -19, 27, -17, 55, -46, -31, -1, 8, -12, 7, -1, 19, 52, -2, 13, 25, 5, 42, 11, 3, -30, -1, -15, -18, 6, 14, -40, -3, 5, -27, -17, -3, 27, -13, 12, 51, 30, -36, -85, 9, -31, 3, 19, 15, 47, -41, -48, -8, 11, 10, 13, 52, 38, -32, -65, -4, 51, 17, -5, 58, -25, -20, -61, -45, -21, 6, 58, 6, 0, -43, -14, -25, 0, -14, 44, 11, 26, -64, 36, -8, 38, -28, 17, 37, 42, 1, 21, -32, -66, 17, 37, 19, -32, -10, -22, 15, -6, -14, 30, 34, -31, 2, 12, 14, 57, 4, -1, 21, 18, -27, 5, -26, -25, 26, 27, -16, 19, 14, 14, 33, 7, -4, 34, -3, 22, -5, 20, -29, 36, 50, -13, 4, -19, 16, -17, 7, 35, -15, 15, -18, 43, -1, 10),
    (-48, 3, 1, 52, -38, 34, -27, 54, 49, 14, -35, 39, -37, 21, 31, 36, -28, 33, -15, -45, 7, -7, -43, -10, -20, -27, -18, 13, 52, -39, 27, 32, -57, 55, -12, -35, 42, -78, -19, -19, -50, 46, 50, 34, -38, 22, -21, -28, -52, -54, -50, -4, -3, 8, 10, -10, -42, -10, 22, -23, 5, -10, -27, 0, -5, -31, 35, 46, 3, -5, 6, -28, -43, 17, -39, 36, -40, -6, 18, 57, 12, -49, -40, 17, -28, 16, 17, 18, 0, 20, 11, -36, -20, -14, -56, -10, 9, -39, -48, -6, -12, -21, 34, 13, -34, 29, -11, -31, 43, -50, -28, 3, 9, 30, 30, 9, -34, 32, 44, -60, 1, -27, 32, -45, 33, -9, 48, -12, -21, 16, 37, 6, -14, 22, -6, 31, 17, 13, -8, -12, 33, 25, -9, -10, 23, 30, -16, -32, 5, -32, 15, 3, 3, -39, 17, 11, -50, 30, -31, 24, -65, -13, -25, -38, 12, 35, 7, 35, 25, -35, -18, 5, -22, -15, 44, 7, -41, -6, -2, -8, 35, -17, 15, -16, 6, 17, -10, 16, 10, 3, -8, -12, 24, -14, 10, -34, -34, -39, 26, -23, -29, 30, 18, -40, 0, -7, 13, 62, -2, -10, -8, 2, 22, -15, 39, 20, -2),
    (67, 4, 9, -21, -20, 2, 31, -4, -38, 12, -5, -2, 24, -11, 27, 7, 8, -18, 19, -37, 54, 42, 31, 28, 25, -1, -14, -25, -10, -39, 4, -18, -73, 39, -23, -13, -29, -9, 29, -36, 59, 40, -8, -33, 34, 22, -8, 28, -2, -27, 32, 26, -6, 5, -24, 22, -52, -12, -16, -31, -12, 27, -9, 18, -52, -6, -12, 36, 34, 38, 33, 34, 10, 41, -20, -67, -19, -37, -23, -13, 38, -39, -7, -7, -41, -36, 19, 55, 25, 30, -37, -13, -4, 29, -16, 55, 3, -28, 24, -48, -26, -34, 28, -36, 25, -30, -12, 27, -32, -13, -59, 4, 92, -12, -19, -58, -26, -20, 33, 3, -118, 17, -15, -2, -25, 36, -8, -43, 28, -14, 24, 27, 14, -7, -40, 44, -18, -62, 9, -44, -22, 9, 0, -36, 4, 23, -42, 16, -26, -21, 27, 19, -4, 26, -29, 17, 48, -33, 24, -28, -7, 40, 0, -19, -1, 53, 10, 5, -1, -45, 34, -10, 16, -53, -36, -51, 44, 20, -24, 16, -42, -30, 23, 12, -4, -2, 6, 12, -67, 2, 23, -20, 24, -13, -62, -48, 1, -8, -15, -103, 41, 42, 21, -12, -29, 18, 9, 5, -22, -37, 3, -2, -54, -53, 26, -10, -6),
    (7, 47, -28, -36, -34, -21, 49, 4, -45, 19, 34, -33, 9, -21, 29, 31, -22, -72, -20, -22, 8, -18, 30, -58, -13, -27, -25, 22, 41, -3, 0, -78, 5, 44, 6, -6, 13, -8, -12, 106, -33, -53, 9, -5, 71, 28, 26, -55, 24, -31, -7, -14, -20, -20, 8, -5, 28, -20, -19, 20, 8, -4, -13, 14, -11, -43, -13, -4, 17, -11, 29, -27, 57, -41, -3, -40, -49, -71, 50, 34, -26, -5, -60, -20, 16, -26, -4, 58, 36, -24, -43, -3, -18, -12, -31, 14, 37, 52, -9, -53, 14, -21, 40, -11, 46, 17, -10, -16, -17, -3, 25, -28, 70, -64, -43, 12, 26, 49, -3, 2, 33, 37, 23, 33, 45, 33, 4, -25, 42, 23, 18, 1, 27, -40, 23, 18, 53, 9, 13, -9, 44, -17, 39, 11, 6, -31, 18, -9, -4, -13, 21, 11, -38, -29, -2, -4, -41, -41, -12, 53, -20, -3, 22, 16, -32, 9, -46, 13, -4, -8, -6, -12, 38, -52, -17, -14, -23, -7, -52, 32, -16, -6, 16, 58, 16, 58, -41, -46, -39, 10, 6, 16, -17, -15, -4, 11, -39, -19, 26, 43, 10, -43, -18, -36, -2, -3, 5, 49, 1, 1, 18, -27, -11, 6, -53, 13, -7),
    (13, -47, -13, -39, 49, 3, -15, -13, -9, 17, -18, -12, 1, -7, -2, -56, -4, -45, 11, 43, -48, -10, 29, -15, 12, -21, 32, -18, 42, -15, 40, -15, 10, 27, -10, 19, -14, -4, -25, -40, -7, -13, -16, 19, -31, -31, -14, 2, -36, -26, 18, 14, -15, -35, 8, -32, 29, 22, -7, 29, -4, 7, 3, -27, 6, 61, -4, 29, -13, -37, 17, -10, -4, -5, 31, -49, -5, -42, -4, -18, 62, -6, -5, 36, 35, -3, -21, 7, 32, -34, -18, -14, 37, -9, -17, -34, -13, 12, -19, 4, -36, 1, 15, 30, -2, -2, 12, -23, -12, 39, 13, -17, 6, 28, 24, -67, 17, 37, 25, -9, 15, -5, 1, 22, -24, 48, 8, 16, -18, -29, -1, -7, 46, 0, -34, -28, 23, 9, 53, 8, -21, 15, 36, -68, -1, 4, -48, -14, 29, -9, -73, -16, -6, 13, -20, -31, -64, -34, 33, -32, -4, 1, -34, -15, -98, 50, -11, 44, -34, -20, 48, -8, 15, 15, -10, 17, 9, -4, -1, 6, -53, -32, 11, -1, -21, 23, -6, 36, -70, 41, -32, 58, -35, -64, -42, -11, -20, 4, -38, -14, 0, 11, -6, -27, -17, -20, 23, 20, -22, 43, 30, 31, -15, 17, -35, 36, -5),
    (-34, -4, -8, -57, -13, -44, -11, -30, -34, -17, -8, 4, -17, -39, -34, -9, 23, 14, 23, 24, -4, 24, 4, -7, 8, -15, 8, -50, -3, -25, -18, 28, -18, -6, -9, 11, 21, 47, -18, 39, -14, 10, 40, -8, 24, 8, 27, -7, 33, -3, 37, -8, 3, -21, -30, 16, -18, -28, -33, -24, -10, -11, 0, -22, 39, 16, 20, 2, 0, 43, 27, 33, 0, -19, -6, -27, -21, -58, 33, 39, -44, 16, 33, -37, 2, -4, -34, 18, -31, -40, -35, 6, -71, -8, -47, 46, 49, 8, 4, 9, -6, -69, -37, 56, -16, -52, -56, -26, -29, 27, 2, 25, 27, -7, 44, -19, -51, 21, -40, 52, 34, 8, -1, -9, 19, -48, 31, -3, 21, 23, -25, 25, -25, -31, 35, 33, 74, 33, 28, -27, -28, 40, 23, 28, -5, 3, -31, 5, 7, -53, 21, -32, 5, 13, -34, -6, -49, -47, 0, 30, -11, -15, -2, -13, -17, -5, -4, -17, 3, 6, -28, 31, -31, -3, 21, 7, 10, -7, -68, 43, 6, -49, 25, 6, 13, 24, 37, 16, -28, 42, 3, 25, 11, -19, -22, 19, -5, 1, 30, 23, 47, 46, -16, -35, 17, -16, 20, -1, 11, 81, 30, -33, -2, 25, 6, 38, -6),
    (11, -22, 7, -16, -20, -60, -8, 11, -5, 26, -26, -18, -21, 31, 48, -13, 44, 46, 53, -25, -29, 8, -19, 3, 36, -9, -30, -33, -6, -12, -5, 30, -26, 9, -18, -2, -12, -45, 13, 4, -1, 29, 1, -2, 44, 27, -26, 42, 40, -19, -20, 26, 35, -12, 16, 2, -4, -35, -36, 13, -12, -14, 3, -18, 44, 0, 55, -12, -1, 9, -20, 7, 35, -7, -12, -3, -49, 22, 26, 18, 52, -32, -24, 33, 11, -24, -24, 50, -18, -21, -19, -35, 69, -8, 18, 13, 73, 37, 58, -22, -18, 28, -9, -4, -10, -30, 33, 39, 15, -2, 35, 8, -19, -6, -47, -53, -11, 16, -42, 31, 9, -13, 29, 67, -6, 32, -19, 47, 15, -6, -58, -7, -40, 49, -18, -34, -19, 39, 35, 25, -10, -18, 10, 73, -10, -14, 22, 20, -46, -46, 2, -32, -15, -39, 38, -24, -15, -16, -18, -3, 22, 19, -17, -4, -39, 9, -16, -38, 3, -1, -14, 18, 21, 58, 17, -24, 24, -23, -18, 27, -28, 35, -16, -43, 25, 42, -16, -2, -16, 21, -22, -1, -16, -5, 28, 15, 24, -3, -36, -25, 9, 31, 17, -24, -4, -29, 22, -8, 3, -2, 38, 10, 27, 42, -17, -1, -5)
  );
  ----------------
  CONSTANT Layer_5_Columns    : NATURAL := 16;
  CONSTANT Layer_5_Rows       : NATURAL := 16;
  CONSTANT Layer_5_Strides    : NATURAL := 2;
  CONSTANT Layer_5_Activation : Activation_T := relu;
  CONSTANT Layer_5_Padding    : Padding_T := same;
  CONSTANT Layer_5_Values     : NATURAL := 24;
  CONSTANT Layer_5_Filter_X   : NATURAL := 3;
  CONSTANT Layer_5_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_5_Filters    : NATURAL := 32;
  CONSTANT Layer_5_Inputs     : NATURAL := 217;
  CONSTANT Layer_5_Out_Offset : INTEGER := 3;
  CONSTANT Layer_5_Offset     : INTEGER := -1;
  CONSTANT Layer_5 : CNN_Weights_T(0 to Layer_5_Filters-1, 0 to Layer_5_Inputs-1) :=
  (
    (0, 48, 0, 20, 11, -38, 32, -8, -71, -24, 16, 17, 7, 23, -18, -23, -59, -15, 6, -11, 24, -31, -9, -13, 10, -19, 4, 15, 27, -34, 40, 23, 1, 38, 18, -17, -62, 33, -51, 12, -52, 13, -4, 64, 30, 45, -29, 8, -1, 21, -13, -27, 52, -31, 42, 21, -35, -9, 19, -27, 3, -11, -40, 13, -22, -21, 34, 11, 5, 26, 10, -21, 41, 23, -21, 19, 26, 0, 52, 38, 17, 31, 31, -2, -17, 13, 12, -30, -48, -9, 21, -9, 2, -14, -5, 28, 26, -14, -22, 21, 54, 21, 59, -47, 8, 30, 0, 4, -47, -39, 7, -1, 15, -24, 27, 32, -8, 82, 26, 28, 32, -16, -8, -7, -4, 6, 65, -1, -11, -11, 23, 35, -50, -55, -29, 3, 17, 4, -4, 10, -59, 40, 23, 32, 16, 24, 23, 9, -15, -19, -2, -8, -27, -21, 12, -8, -52, -15, -11, -34, -15, -19, 21, 13, -12, 37, 10, 5, 44, -4, 51, -44, 24, -35, 27, -35, -8, 62, 21, 6, -66, -36, -10, -22, 26, -23, 24, 32, 3, 14, -17, 50, 1, 44, 39, -40, 6, -29, 40, -56, -26, 40, 8, -37, -8, 0, 26, 12, -1, -23, 1, 18, -48, 15, 23, 24, -2),
    (-15, -15, -42, 39, -22, 40, 20, -10, -21, 26, -11, -13, -28, -34, 26, 7, 32, -12, 10, -10, -49, -11, 41, 11, -17, 5, -22, 60, -33, 38, -28, -16, 19, 27, -39, 8, -17, 52, 16, 1, 8, 3, 60, -54, -34, -43, -31, -10, -5, -3, -8, 33, -34, -4, -31, 23, 6, -8, -35, 11, 11, 7, 6, 39, 15, -25, 35, -34, -11, -41, -40, 16, 9, -17, -58, 57, -5, 28, 0, -8, -13, 37, -16, -13, 27, 6, -3, 1, 2, -6, 57, -68, -39, -67, 16, 34, -27, 20, -28, 54, -45, 45, -30, 10, 39, -7, -42, 14, 55, 25, 40, -1, 9, -33, 45, -10, -10, -35, 22, -21, -1, -47, 29, 47, 47, -21, 25, 39, 5, -29, -27, -8, 56, 0, 45, 13, 17, -27, 61, -46, 0, 5, -13, 17, 29, 34, -19, 16, -10, -29, -16, 7, -33, -51, -35, 11, 14, 36, -17, -15, 13, -9, 48, -66, 17, -61, -17, 5, -14, -37, 4, 28, 28, 10, -3, -27, 7, -12, -65, 9, -6, 45, -9, 12, -2, -13, 35, -44, 27, -2, -7, -3, 9, -22, 26, -39, 33, 36, 12, -29, -41, -24, 17, 37, -31, -25, 38, -15, 21, -12, 7, 8, -1, 7, 31, 30, 5),
    (-9, -3, 14, 6, -8, -27, 20, -29, 15, 12, 9, 4, 16, 9, -39, -2, 25, -8, -22, -41, 22, 11, -1, -3, -62, -38, 9, 25, -2, 25, -6, -37, -10, 7, -30, 1, -19, -10, -19, -29, 7, -2, -26, -38, 28, 38, -8, -13, -51, -29, 20, -12, 3, 18, -17, -33, -54, 12, -30, -18, -37, -43, 19, -39, 19, -37, 21, -19, -30, 21, 1, -13, 33, 43, 69, -31, -10, -24, 12, 45, -8, 42, 27, 38, 26, 36, 20, -43, 11, -17, -22, 50, 43, 45, 36, 41, 16, 62, 65, 23, 9, -41, 4, 37, -50, 56, 15, 4, 48, 10, 13, -33, 55, -30, -5, 45, 37, 27, 12, 32, 8, 24, 4, -29, -14, -16, 18, -8, -37, 22, -2, 4, 8, -31, 4, -4, 50, -38, 38, -10, 23, 59, 27, 3, 19, -18, -23, -15, 29, -28, -3, -5, 3, 34, -42, 25, -32, -16, 12, -27, 9, 0, 27, 34, 20, 7, -30, 10, 18, 8, -26, -17, -11, 27, 5, -8, -33, 23, 2, -2, 12, 2, 29, -27, -7, -9, 0, 2, -32, 44, -5, -6, 17, -6, -4, 23, -7, 0, 30, -11, -20, 15, -19, -16, 8, -23, 11, 46, -18, 32, 14, -40, -20, -24, -43, 6, -6),
    (-46, -5, -62, 20, 44, -1, 42, 22, 13, -29, -52, -1, 8, 2, -10, -14, -27, 11, -6, 55, 56, 36, -2, 33, -30, -42, -21, 23, 19, -30, -33, -20, -34, -37, -62, -42, 30, -26, 2, 5, -46, -46, -28, 34, -30, 1, -37, -11, -29, -42, -23, 2, -13, -31, -65, -40, 43, -50, -79, 12, 28, -16, -10, 4, -23, -5, -19, -22, 17, 22, -64, -25, 29, 17, 24, -24, 34, -29, 23, -26, -19, 38, 11, 15, 11, 49, -44, -50, 8, 1, -52, 37, -3, 14, 39, -21, 28, -4, 25, -3, 32, 31, 40, 40, 10, 35, -24, -34, 74, 10, -50, -26, -2, -23, 24, 41, -16, 42, 35, 3, -23, 2, 28, 10, -27, -18, 20, 2, 27, 41, -28, -39, -12, -29, -6, 4, -15, -53, -34, 25, 18, -16, 14, -3, 4, -10, 3, -2, 35, 18, 0, -18, 4, -27, 45, 22, 8, 34, -37, -19, -5, 31, -16, -3, -42, -21, 5, 10, 46, -15, 28, -12, -19, 43, 58, 0, 4, 23, -10, -22, 21, 23, -23, 27, 33, 26, 8, 28, -50, 35, 7, 28, -12, -9, 49, -66, -33, 22, 0, -6, 8, 20, 23, 0, 6, 3, -40, 23, -22, -13, -14, 25, -18, 8, -5, 20, 6),
    (3, 37, 3, 22, 50, 31, 49, -13, 11, -3, -31, 8, -19, 16, -17, 14, 35, 30, -4, 59, 25, 45, -2, -9, 20, 44, 15, -5, 27, -33, 23, -27, 30, -3, -37, 14, 2, 0, 30, -40, 25, -15, -8, 53, 58, 51, -7, 17, -8, 35, 9, 12, -6, 16, 9, -14, -36, -30, -11, 17, 5, -3, -13, 5, 30, -16, -23, 13, 31, 23, 6, 10, 1, -14, -1, 7, 79, -2, 49, -12, -6, 29, -21, 16, -40, -20, -21, 18, 32, 22, -24, 77, 49, 36, 17, 38, -24, 53, -14, -54, 93, -7, 17, -43, -9, 20, -20, -14, -31, -12, -12, 8, -8, -18, -64, 77, 40, 64, 41, 61, 4, 50, -16, 8, 62, -34, -17, -30, 7, 23, -43, -43, 7, 28, -30, 19, 10, -32, -69, 25, -15, 33, 17, 70, -17, -2, -15, -32, 57, -33, 17, 19, -25, 0, -34, 25, 13, 10, -27, -12, 11, 17, 5, 35, 41, 16, 26, 36, 19, 24, 10, -37, 45, -22, 18, -18, 2, -34, -15, -6, 9, -10, -37, 10, -16, -12, -27, 32, 49, 8, 11, 62, 6, 23, -31, -40, -26, -3, -32, 27, -14, -42, -36, -23, -27, 18, 10, -16, 12, -1, -54, -10, -2, -34, 14, 27, -7),
    (47, -27, -28, -4, 26, -9, 8, -40, -70, 13, -73, 14, 39, -37, -19, -59, -1, -25, 24, -13, 3, -22, 23, 26, 45, 13, 8, 17, -5, -35, 8, 10, -54, -32, -33, 8, -22, -39, -38, -11, 36, 13, -61, -16, 34, 5, -25, -14, 42, -27, -22, -6, 0, -20, 26, -63, 19, 12, 17, 16, -10, 0, -11, -21, 19, -18, -46, -12, -32, 43, 31, 16, 31, 3, 0, 26, 8, -36, 7, -35, 12, -1, -48, -42, -38, 3, -19, -46, -5, -9, -5, 4, -10, 32, 22, 31, 1, 3, -16, -10, 43, 5, 60, -29, 25, 16, 32, 6, -3, -21, -62, -21, 24, 8, -63, -6, 25, 46, 5, 43, -1, -10, -26, 0, -13, -5, 23, -34, -30, 24, 1, -35, 6, 21, -32, -39, 4, -23, -5, 31, -2, 29, 29, 18, 0, -32, 3, 11, 15, 14, 27, 23, 7, 19, 36, -38, 6, 37, -56, -28, 27, 30, 26, -10, -13, 19, 5, 11, 21, 32, 13, 14, 53, -17, 42, 17, -26, 7, 30, -48, 11, 38, -33, 10, -30, 22, -8, 22, -35, 21, 58, 45, 8, -27, 1, -14, 57, -29, 29, 9, -21, 21, 2, 8, -13, -19, 3, -5, 33, 11, 36, 12, -4, 42, 8, 22, -3),
    (25, 25, 33, -16, 59, 19, 3, -18, 60, 7, 4, 36, 7, -2, -23, -45, -16, 12, -11, 35, -7, 42, -7, 20, -17, 19, -12, -12, 63, -37, 33, 34, 21, 29, -18, 16, 12, 15, -45, 12, 14, 9, 0, 4, -20, 38, 5, 5, -11, 21, 33, -15, 50, -26, 42, 43, -9, 1, -21, 1, -2, 30, -39, -8, -9, -15, -16, 24, 16, -20, -12, -15, -10, -22, 16, -5, 1, 6, 43, -26, 70, -71, -38, -27, 41, -52, -27, -57, -35, 9, -39, -22, -43, -48, -33, 46, -41, -6, 20, 14, 1, -12, 26, 8, 8, -16, -14, -17, 14, -61, 18, 6, -26, -48, 4, -59, -40, -23, -44, -41, -54, 7, -52, 7, -11, -2, -20, -21, 55, -55, -55, 18, 24, -37, -3, -42, 14, 2, 41, -53, 2, 2, -15, -26, 2, -13, -43, 21, -34, -32, -19, -45, -29, -3, 9, -40, -18, -9, -28, -39, -4, -30, -32, -9, -8, 37, -16, 6, -45, 14, -22, 23, -1, 6, -8, -2, 32, 19, 18, 34, -37, -24, 34, -35, 46, 9, -10, -15, 5, 35, 2, 46, -1, 5, -20, 62, -14, 8, -15, -78, 18, -5, 27, 35, 0, 10, -5, -1, 37, 3, 47, -59, 14, 37, 39, -1, 2),
    (-13, -39, -12, 6, -34, -16, 40, 14, -53, -7, 40, 8, -24, 18, 34, -32, -7, 1, -23, 0, 29, 50, -26, -35, 22, -18, 4, 26, -4, -26, 47, 18, -27, 36, 17, 35, -48, -11, -15, -2, -38, -48, -3, 35, 56, -21, -4, 9, 3, -13, -5, -2, 7, -26, 8, 11, -5, -29, 15, 6, -20, -13, 21, -35, -22, -16, -6, 50, 1, 1, 14, 21, -36, -4, -29, 56, -4, -35, 12, -11, 23, 16, 15, -14, -61, 63, -49, -39, 25, 20, -43, -47, -29, 20, -7, -2, -27, -5, -16, 73, 5, -7, 23, 11, -26, 22, 29, -65, -44, -12, 8, -65, -13, 40, -49, 19, 20, 8, -49, -33, -31, -28, -6, 17, 1, -15, 33, 26, -22, 19, -21, -40, -47, 11, -8, -55, -49, -38, -38, -20, -34, 0, -7, -39, -15, 44, 16, -3, 8, -36, 75, 22, -34, 48, -5, -37, -15, 47, -39, 6, -15, -20, -7, 24, 8, 38, 4, 50, -39, -36, 34, 16, 20, -4, 79, 4, 15, 53, 25, -24, 27, 29, 14, -60, -31, 5, 2, 20, 19, 28, 4, 66, -24, 18, 11, 14, 9, -23, 48, -43, -17, -10, -21, -42, 24, 39, -1, -10, 39, -29, -16, -11, 34, 16, -19, -25, -2),
    (-30, -10, 24, -1, -8, 23, 9, 1, 7, 16, 0, 4, 41, 6, 3, -11, -3, 45, -7, -16, -45, -12, -16, -20, -21, 7, 43, 43, -16, -42, 39, -37, 47, 44, 32, -9, 31, 6, -47, 1, -17, 18, -20, 19, 4, 14, -2, -35, 1, -3, -4, 65, 25, -14, 17, -29, 28, 6, 9, 9, -18, -13, -22, -23, 20, 20, 20, 30, -9, 25, -5, 24, 5, -12, 60, -60, 18, 11, -29, 9, 27, 48, 68, 36, 21, 0, -1, -31, 26, 55, 45, 3, 7, -34, -14, 4, 56, 49, 71, -39, -5, -35, -16, -7, 7, 25, 24, 3, 35, 25, 16, -33, -4, -4, 22, 12, 33, -21, -8, 26, 15, 37, 29, 11, 20, -33, 12, 15, 51, 23, 62, 10, 5, -37, -2, -31, -16, -11, 1, -16, 54, -19, -37, 21, 40, 56, 57, -38, 11, 17, -15, -4, 29, -20, 56, 30, 21, -38, -6, -29, -30, -10, -10, 6, 17, -36, -33, -34, -3, 10, 14, -35, -20, -37, 7, -7, 49, -29, 9, 40, 12, -57, 20, -20, 9, -32, 32, -13, 28, -37, -58, -33, -22, 18, -10, -9, -43, -3, -53, 10, 17, -63, 30, 39, -8, -31, -21, 17, -22, -35, -8, 11, -2, -24, 17, -35, -6),
    (-11, 8, 15, 14, 34, 23, -57, 11, -14, 7, 16, 0, -17, 42, -7, -23, 20, 24, 8, -35, -19, -11, -7, -39, 28, 5, 4, 2, 39, -23, -13, 8, -58, 29, -29, 14, 18, 56, 34, -30, 17, -6, 43, -5, 23, 35, 15, 6, -3, -18, -15, -40, 22, -32, -9, -41, 1, 43, -17, -4, 4, 30, 9, -7, -43, -24, 26, 3, 4, 45, -1, -39, -24, -7, -52, -37, 59, -16, -3, 13, -21, 22, -6, 11, -41, 36, 23, -17, -18, 15, 25, -28, 7, 41, -34, -30, 0, -33, -21, -39, 33, -32, 73, -3, -33, 57, 3, 41, -40, 36, 30, -2, 3, 16, -15, 22, 29, 77, -13, -5, 23, -19, 15, -29, 70, 26, 42, 27, -32, 66, 10, 7, -4, 26, 26, -8, 26, 31, 1, 18, -38, 53, -15, 26, -32, -5, -36, -2, 54, 20, -16, 2, 19, 41, 15, -4, -5, -4, -8, -7, -3, 16, -3, -2, 3, 23, -19, -15, -24, -34, -43, -40, 20, 39, 0, -6, -43, 43, -20, 10, -31, 33, -12, 20, -15, 7, 35, -11, -26, 38, -42, 20, -21, -14, 14, -45, 20, 43, 9, 2, 2, 9, 40, -21, 19, 33, -9, -26, -16, -6, -64, 22, -31, 61, 5, -21, -12),
    (50, 1, -13, -29, 10, -34, 8, -23, 32, 9, 18, -31, 20, -49, -40, 20, 2, -52, -46, 63, 3, 58, 29, 33, 8, -4, 23, -22, 7, 10, 31, -23, 21, 20, 58, -41, -8, -13, -24, 22, 7, 28, -20, 51, -25, 51, -24, 24, 25, 32, 32, -10, 15, 8, 11, 39, -21, 40, -25, 10, -39, -10, 13, 20, 30, 21, 29, 46, 14, 38, -20, 20, 35, 3, 13, -33, 17, -24, 37, 41, 7, -8, 42, -21, 17, -22, 19, 8, 16, 22, -29, 35, 35, 13, 21, 12, 57, 27, 45, -15, -14, -30, 57, 10, 26, 19, 71, -45, -8, -26, -18, -21, -31, 5, -35, 79, -16, 68, 26, 61, 34, 38, 61, -15, -26, -4, 31, -5, 12, 5, -2, -38, 6, -16, -25, 30, -6, 42, -8, 33, -15, 26, -2, 33, -17, -30, 20, -15, 21, -33, -7, -6, 38, 31, 54, 0, 14, -30, 9, 42, -9, 27, -18, 6, 19, 9, -3, 18, 19, -3, -2, -22, -5, 11, 30, 22, 34, -2, 34, 4, 23, -7, 4, -22, -25, 18, -8, 39, -11, 28, -9, 25, 25, -19, 40, -6, -56, 43, 36, 0, 51, 7, 17, -14, -28, -54, -33, 0, 17, 20, -41, 12, -5, -7, 25, 9, -4),
    (36, -38, 30, 46, 10, 0, 10, -13, 13, -13, 22, 19, -18, 22, -40, -9, -36, -19, -13, -16, -15, 24, 67, -18, 42, 18, -34, -8, -56, 8, -9, 21, 57, -9, 18, 7, 14, -12, -41, 36, 2, 16, -19, -16, 39, 25, 74, 27, 9, -5, -8, -27, -12, 2, -6, 46, 22, -2, 47, 12, 2, 50, -3, 24, 23, 56, 36, -23, 29, 18, -10, -18, -10, -25, -10, -44, -28, -17, 35, -14, 17, 26, 32, -19, -73, -68, -30, 33, -4, -8, 3, -17, 15, 68, 28, 54, 52, -10, -51, 22, 0, 11, 42, 13, 52, -5, -5, -8, -34, 0, -31, 64, -35, 33, 20, -1, -10, -8, -8, 25, 26, 21, -16, 42, -25, 23, -16, 2, 30, -18, 20, 1, -40, 23, 23, 59, -15, 39, -4, -9, -14, -2, -15, 10, 7, -18, -45, 16, -6, -48, -7, 21, 29, 14, 27, -46, -26, -12, -52, 8, -12, 41, 13, -32, -10, 19, 31, 39, 23, 23, -34, 32, -5, 11, 21, 6, 16, -24, 1, -34, -30, 6, -31, 4, -44, 59, 15, -49, 1, 24, 31, 2, -26, 24, -10, 35, -14, -7, 14, -20, -1, -44, 0, 15, -37, 9, -2, -2, -64, 13, -1, -16, 15, -45, -47, 36, -2),
    (-18, -10, -21, -3, 2, -2, 56, 3, -17, 36, 38, -11, -36, 35, -24, -14, 19, 45, -39, -8, 2, 6, 28, 10, -47, 10, 4, -2, -9, -24, 32, -32, -43, 9, 15, -81, -5, 23, -34, 4, -6, 22, -15, -31, -35, -14, -50, 17, -14, -1, 15, 42, 5, -22, -10, -34, -21, 23, 7, 2, -46, 4, 6, -38, -34, 31, 2, -61, -58, -35, 15, 13, -9, 19, 40, -30, 45, -7, 23, 20, -11, -13, -28, 9, -31, -15, 2, 37, 39, 11, -36, -5, 21, 39, -30, 53, -21, 25, 60, -24, 26, -16, 13, 22, 7, 36, 3, -12, -50, 21, -9, -25, 40, 34, 4, -29, -34, 2, -1, 8, -61, -17, 44, 23, -25, -13, -12, -39, -16, -5, -28, -38, -26, 33, -28, -16, -13, 4, 22, -16, -34, -37, -41, -9, 25, 27, -5, -3, 31, 5, -21, 42, 0, 11, -21, -38, -19, 7, -19, -30, 11, 15, 14, 15, 35, 33, -33, 51, -22, 0, 55, -1, 7, -9, -25, -36, -56, -2, 23, -2, -20, -23, -18, -2, 4, 31, -10, 18, 16, 6, -3, 31, -49, -18, 54, 6, 3, -12, 27, -13, -33, 23, -12, -25, -27, -3, 19, 33, 22, -22, 31, -20, 13, 8, 26, 49, 0),
    (-32, -20, -23, -14, 12, -33, -32, 37, 51, -15, 15, 21, 41, -38, 7, 3, -16, 43, -24, 5, 24, -17, 29, -2, 20, -42, -24, -32, -1, -7, -44, 14, 51, -26, -1, 23, 73, -3, -22, 18, 3, 37, -38, -15, -23, -43, -17, -16, 16, -74, -45, 10, -42, -16, -33, -13, 26, -30, -23, -32, -1, -64, -43, -14, -26, -47, -35, 3, -12, -38, -53, -30, 31, -13, -7, -31, -5, -35, -16, -12, 10, -48, 0, 28, 60, 18, 5, 34, 3, -6, 33, 19, -1, -1, 34, -36, -22, 18, -1, -52, -45, 28, -27, -28, 11, -36, 15, -39, 54, -33, -31, 6, 19, 16, -18, 21, 1, -19, -36, -37, -23, -2, -39, -8, -63, -32, -30, -11, 35, -60, -53, -39, 47, 0, -9, 21, -39, 0, -40, 35, 35, -27, -66, -30, 20, 25, -12, 5, -59, 7, -13, 23, 46, 33, -1, 26, 61, 10, 27, -26, 32, -20, 17, 8, 3, 27, 27, -24, -24, -20, 7, -2, -54, -39, -8, -17, 64, -11, 23, 18, 91, -9, -6, 20, 11, -42, -30, 32, 33, 65, 53, 13, 25, -36, 1, -33, -18, 14, -16, -32, 20, -2, 23, -28, 20, -4, -13, -19, 1, 11, -48, 38, 27, 40, -11, 4, -1),
    (22, 3, 15, -9, 9, 15, 37, 19, 4, 21, -5, 19, -62, -3, 56, 31, 6, -29, 7, 10, -2, -13, -32, 28, 16, 53, 55, -38, -26, 33, 31, 50, 3, 51, 38, 41, -18, 28, 28, 9, 27, -2, 18, 38, 19, -8, 0, 18, -2, 21, 56, 2, -29, -33, 9, 12, 27, -6, 49, 42, 25, -13, 21, 20, 36, 14, 3, -1, 19, 14, 20, 22, -2, 6, -11, -4, -25, 0, 26, -1, 25, -46, 6, 11, -58, -11, 20, -15, -8, -39, -11, -9, -10, -46, -39, 18, -16, -7, 17, -24, -95, 3, -5, 61, 24, -29, 43, 30, -63, -39, -15, 13, -1, 8, -21, -45, 8, -63, -10, -23, 20, -15, -19, -9, -74, 45, -6, 50, -5, -47, -3, 29, -21, -13, -21, -2, -14, 1, 26, -38, -40, -42, 17, 13, -8, -11, -56, 43, -2, -20, -12, -45, -21, -34, -22, -18, -52, 2, -25, 6, 12, -1, -1, -27, 25, 13, 4, -23, 18, -7, -21, 45, -34, 14, -1, 35, -25, -12, -29, -10, -73, 19, -20, -28, -42, -26, -14, -64, 2, -72, -40, -28, -44, -31, -56, 32, -16, 3, -25, 47, -19, -18, -34, -41, 18, 32, -3, -21, -32, -20, -20, -38, -40, -34, -28, -44, -11),
    (-3, -5, 36, 24, 32, -8, 34, -38, -11, -8, -42, -23, 2, -44, -37, -12, 7, 17, 7, 38, 3, 40, 49, 36, 40, 28, 18, -9, -21, -30, 29, 19, -50, 63, -18, 20, -24, -24, -33, -13, 8, -16, -2, -12, -24, -4, 11, 32, -19, -19, -41, 45, 13, 0, -3, -33, -35, 35, 22, 7, -19, -20, 24, 19, 3, -17, 32, 8, -9, -13, 23, -2, -15, 16, 44, 4, 18, -12, 23, -28, -8, -18, -32, 6, -9, -30, -25, 23, 10, -21, 19, -9, -7, 12, 40, -6, -17, 11, -4, -24, -14, -38, 42, -11, -14, 24, -9, 24, -2, -64, -46, 47, -47, -19, 0, -26, -25, 15, 73, 16, 6, -31, 3, 34, 12, -32, 38, 0, -31, 37, -14, -12, -13, 5, -2, 29, 21, 17, 42, 0, -2, -16, 57, 18, -19, -14, 21, -25, -19, -39, 47, -10, -2, 57, 15, 7, -34, -17, -22, 17, -26, 1, -6, 26, -1, 23, 54, 12, 3, -32, 15, -14, -19, 35, 60, 6, -58, 56, -14, 7, -8, -51, -22, 42, 4, -45, 32, -2, -60, -6, 16, 18, -35, 17, 0, 3, -13, 3, 7, -8, -20, -23, -15, -34, -37, 20, -5, 36, 15, 3, 22, -26, -6, 20, 53, 35, -2),
    (48, -13, 41, -59, -15, 27, -5, 4, -17, 33, 16, 49, 37, -10, 26, 47, 7, 4, -29, 24, -1, -28, -64, -35, 9, -13, 13, -78, 52, 5, 7, -26, 28, -22, 12, 51, 47, -17, 28, 15, -5, 22, 16, -9, -4, 16, -29, -43, 9, 2, 1, -21, 16, 8, -3, -14, 25, 14, 25, 35, 7, -25, 23, 32, 10, -36, 2, -15, 33, -8, 30, -13, 19, -10, 42, -47, 25, -34, 23, -17, 0, -14, -40, 49, -7, -55, 12, 33, 29, -15, 25, 5, 25, 39, 19, -10, 38, 21, 32, -91, 49, -20, 57, -35, 17, 66, 3, 40, -22, -32, 47, -6, -27, -17, 4, 16, 14, 52, 25, -18, -6, -19, 46, -103, 24, 24, -18, -13, 37, 45, 35, 31, -6, -25, 8, 10, 4, -37, 1, 25, 9, -3, 16, -15, -28, 32, -8, 3, 22, -10, -3, 17, -16, -7, 13, -9, -49, -10, 5, -2, -30, 8, -38, 41, -14, 5, -14, 12, 31, 3, -26, -62, -3, -8, -9, -17, 5, 25, -3, -8, -63, -52, 20, -36, 25, -38, -42, -10, -62, 12, 20, 28, 33, -19, -45, -15, -46, -2, -40, -57, -18, 46, -40, -32, -23, -42, -32, 0, -4, -70, 2, -36, -65, 38, 25, 21, -7),
    (27, 2, 11, -21, -12, -14, 9, 8, -3, 24, -16, 11, 14, -31, 25, -49, 6, 25, 6, 16, -31, 32, 68, 18, -39, -11, 44, -41, 26, -5, 3, -8, -3, 68, 25, 31, 3, 14, 5, -10, -27, -55, 7, 39, 12, -1, 60, 8, -40, 3, 28, -52, 22, -14, 12, 29, -31, 45, -20, 17, 21, -8, 3, 4, -23, -17, 20, 11, 26, 29, 18, -16, 27, -55, -24, -46, 24, 33, 11, -70, -91, 55, -41, -4, -7, -8, 18, -59, -28, -43, -12, 18, -5, 24, 72, 78, -24, -24, 23, -47, 16, 49, 8, -22, -1, 90, 9, -21, 20, -26, -33, -2, -31, -63, -4, 22, -43, 15, 75, 55, -45, 17, 35, -13, -15, 46, 10, -22, 16, 45, 8, 8, 32, -4, 11, 1, -36, -25, -42, 17, -55, 34, 12, 37, -1, -38, -13, -3, 57, 29, -33, -46, -13, 31, -32, 1, -40, -40, -5, -15, 15, -12, -31, 14, 30, 5, -12, 47, -5, -3, 13, 14, 15, 14, 10, -44, -6, 54, 14, 20, -14, 2, 24, 0, -21, 6, -5, 10, 1, -8, 59, 34, -25, 8, 12, 4, -5, 34, -26, 2, 12, -11, -5, -8, 45, -28, 10, 43, -21, -19, 20, 3, -16, 20, 27, -7, -8),
    (-35, 1, -15, 30, 11, -36, -7, -12, -18, 13, -36, -50, -12, -19, 1, 35, -13, -24, -37, -12, -38, -15, 11, 17, -39, -53, -5, -20, 18, -24, 22, 5, 1, -14, 42, -59, -46, 8, -56, -8, -22, 1, -34, -33, -30, 10, 36, 17, -51, -14, -30, -27, -11, -37, 13, -14, 21, 8, 43, 7, -38, -18, -9, 2, -4, 29, 6, -42, -68, -3, 12, 5, -31, -12, -31, 21, 22, 27, -10, 28, -23, 23, -6, -45, -81, -36, -52, -4, -18, 2, -11, -16, -7, -14, 21, 27, -32, 10, -40, 4, -26, -28, 23, 29, 19, -18, 18, -52, -35, 35, -32, 0, -22, 50, 49, -59, -29, 4, -21, 9, 11, 19, -41, 35, 15, 20, 13, 62, 56, 19, -2, 1, -19, 11, -40, 4, 31, 55, 20, -64, -39, -24, -33, 6, -30, -17, -17, -14, 16, 34, -1, -3, 20, 21, -29, -48, -18, 3, -48, 41, 17, 19, 28, -19, -9, 4, -21, -14, 15, -18, -26, 31, -20, 14, 20, 47, -4, -21, 16, -36, -77, 46, 2, 34, -9, 51, 45, -59, -11, -12, -14, -24, 2, 37, -8, 29, 56, 5, 24, 36, 1, -3, 52, 1, -49, 44, 42, -15, -15, 58, 13, 1, 3, -11, -31, 7, 18),
    (-8, -24, 4, -11, 28, -27, 7, -44, -35, 5, -15, 54, 19, -30, 17, -2, 4, -41, 10, 19, -9, -5, 4, 52, -23, 32, 33, -19, 28, -14, -9, -28, -47, 6, -15, 6, 4, -19, 51, -2, 2, -64, 44, 0, 29, 13, 33, 14, 32, -4, -8, 15, 21, -16, 19, -16, -4, -15, -48, 22, -25, -1, 39, -26, -1, -5, -5, -19, 51, -4, -2, 7, -3, -47, -30, -40, -15, 8, 31, 8, -22, 25, -9, -4, 27, -33, -4, -30, 8, -23, 25, -2, 28, -12, 16, 23, -36, -34, 19, 10, 24, 33, 45, -21, -50, 0, -43, 56, 27, 12, 25, -12, 32, -75, 59, 9, 9, 0, 45, 47, 20, -1, 14, -7, 0, 12, 18, -15, -5, -7, -42, -7, -24, -3, 21, 19, 39, -30, 5, -39, 8, 21, 35, -42, 18, -51, -20, -58, -37, 25, 17, -19, -9, 40, 16, 29, -39, -32, 0, -12, -10, -19, 3, 21, -23, 11, -4, 3, 20, -33, -13, -4, 26, -23, 10, 23, -35, 43, -36, 41, 12, -36, -9, -38, -19, -16, 0, -3, -29, 14, 9, 32, 21, -17, 11, -2, 1, 14, 2, 45, 12, 4, 18, 25, 6, -18, -15, -4, 34, -11, 27, 24, -24, -2, 37, -10, -12),
    (-25, 1, -14, 3, -25, -33, -25, -28, -24, 9, 21, 1, 43, 7, 34, -45, 50, -8, -1, 10, 28, 18, 34, 15, -11, -37, -19, -2, 2, -20, -45, -41, -16, 7, 1, -33, 54, 18, 38, -34, 54, -19, -7, -6, 59, 31, 1, -5, -18, -44, 18, 9, -3, -32, -30, -24, 17, -5, -13, 17, -31, -2, 7, -1, 24, 3, -29, 33, 57, -8, -23, -33, 24, 30, 14, -33, 20, 26, -19, -37, -5, 21, 34, 53, -34, 54, -35, -29, -31, 12, -13, 44, -20, 18, 37, -38, 38, 44, -5, -86, 23, 7, -10, 30, 10, 44, 46, -6, -12, 25, 0, 4, 47, -21, -3, 32, 35, 13, -6, 30, 6, 32, 17, -37, -9, 5, 48, 15, -21, 54, 26, -24, -39, -32, -28, -2, -16, 22, 14, 27, 14, 31, -7, 30, 8, 0, 19, -46, 0, 8, -20, -15, -15, -4, -6, 14, 7, 21, 3, 13, -44, 9, -22, 5, -18, 13, 23, 6, 8, -25, 44, -16, 33, 13, 7, -15, 0, 47, 3, 39, 57, -53, 12, 0, 5, -3, -27, -3, -12, 12, -11, -5, 37, 7, 56, -7, -21, 14, 42, -11, -7, 32, -13, 22, 49, -34, -44, 9, -22, -33, -1, -4, -13, -11, -3, 36, -8),
    (-31, 26, 39, -58, -27, 18, 12, -41, -5, 21, -16, -30, 8, -9, -40, -6, -15, -30, 53, 5, -7, 12, -10, -20, -75, -26, 10, 10, 8, -2, -5, -46, 22, -29, -32, -5, -25, -37, -52, 43, -27, 28, 16, -13, 30, -52, 54, -3, -78, -33, 2, -10, -51, -28, -34, -59, 43, -59, -49, 15, -26, -34, -22, 41, 27, -2, -13, -31, 40, -21, 41, -2, 10, 18, 39, 1, -24, 7, -2, 0, -15, -17, 29, -22, 23, -24, -57, 21, -21, -4, -21, 32, 39, -12, 17, -2, -57, 47, -2, -8, -46, 23, 11, -29, 48, 3, -44, 3, -8, -70, -28, 69, 32, 5, 9, -13, 39, -6, -12, 31, -67, 3, 6, -6, -23, 6, 0, 16, 43, -1, -3, 37, -20, -41, -31, 55, 14, 7, 17, -29, 15, -5, 13, -31, 10, -31, 40, -63, -1, -18, 12, 29, -36, 33, 19, 43, -40, -49, 16, -3, 16, 19, 4, -12, 30, 20, 6, 17, -5, 15, 28, 9, -45, 50, 12, 20, -25, -10, 19, 12, 31, -53, -41, 38, 50, -44, -37, 13, 0, -11, -27, 45, 17, 21, 19, 15, -45, -3, -16, -11, -1, 3, -29, 30, 7, -43, -12, 10, 32, 33, -34, 17, -16, 6, -16, 2, 3),
    (-44, -6, 7, -1, 23, 27, -12, -23, -36, 44, -12, -24, 5, -27, 4, 15, 17, 11, -12, 42, -12, 20, -29, 3, 1, -50, -16, -4, -15, 38, -17, -35, -7, 14, -72, -2, 28, -2, 12, -76, 9, -28, -1, -3, -17, 40, -34, 9, -64, 3, -18, 28, -21, 19, -30, -56, -6, 15, -19, 21, -25, 8, -27, -13, -1, -9, -25, -14, -34, 8, 3, 1, -9, -15, 34, 31, -23, 40, -67, -21, -29, 37, 9, 31, -18, 15, 32, 13, 9, 6, -20, 9, 5, 20, 7, -38, 0, -29, -6, -35, -19, 13, -16, -32, -6, 38, 12, 22, 2, -13, 41, -21, 69, 21, -15, -29, 8, -11, -31, -34, 11, -8, -20, 18, -10, 10, 52, -40, -20, 21, -18, 27, -13, -33, -15, -53, 24, 6, 15, 13, -22, 14, -24, 33, 19, 28, -15, 0, -26, 8, 14, 18, -49, 30, 27, -31, -9, -16, 9, -67, 23, -12, -7, -7, 6, 1, -25, 6, 35, -23, -1, -32, -59, 19, 31, -4, 9, -14, 58, 19, 28, -41, 32, -51, 48, 50, 20, 7, -17, -16, -52, -13, 20, -24, -29, 3, 15, -14, -3, 29, -47, -2, 35, 40, -15, 3, 16, -53, 34, 53, 10, -9, 22, -17, -3, 42, -4),
    (-2, 27, -5, 30, 24, -7, -27, 2, -29, 42, -10, -4, 17, 13, 11, 3, 38, -26, 31, 36, 32, 28, 21, 32, 48, -17, 21, -32, 38, 8, -31, -3, -62, 9, -18, 21, -4, 24, -27, -45, 15, -56, -13, 43, 5, 50, 28, -7, 14, -27, 29, -16, 29, -1, 14, 36, -38, -5, 36, -26, 29, -34, 1, 19, 2, -45, 3, -19, -22, 12, 15, -21, -23, -15, 2, -25, 34, 28, -10, -25, 5, 41, -1, -25, 14, -1, 3, -7, -14, -19, -23, 61, 20, 58, 26, 0, -16, -2, 53, -43, 38, 31, 37, 2, 6, 50, -61, 13, 30, -6, 17, -27, 4, -11, -45, 62, -44, 35, -16, -28, -60, 1, 42, -3, -5, -25, -17, 13, -30, 24, -51, -6, 34, -28, 15, 17, -58, -25, -56, 23, -73, -4, -67, -29, -27, -12, 32, -36, 37, 14, -10, -26, 37, 34, -28, 23, -8, 4, 33, 46, 28, 7, -9, 8, 16, 29, 38, 36, -40, 14, 30, -27, 43, 38, 34, -30, 53, 37, -28, -16, 0, 33, -13, -46, 29, 9, -37, -10, -6, 6, 47, -40, -34, 17, -39, -13, -13, -26, -20, 17, 37, 3, -8, -53, 0, -8, -47, -28, -25, -27, -51, 38, -26, -17, -6, -66, -9),
    (-57, -20, -5, -12, 13, -20, 7, -39, 5, 9, 24, -58, 68, 5, -31, -5, -15, 19, 19, -25, -28, -49, 10, 10, -61, 28, -20, -29, 2, -13, -15, -57, 9, -53, -9, -15, 10, -44, -12, 16, 22, 13, -5, -41, 26, 19, -24, 28, -10, 31, 6, -30, -19, 19, 15, -67, -29, -18, -19, -43, 11, -2, 11, -35, -47, -17, 40, -7, 22, -48, 45, -62, -30, 6, -44, 22, 6, -9, -35, -5, 37, -27, -41, 22, 73, -43, 43, -2, 21, -38, 6, -16, 14, 20, 16, -12, -35, -28, -13, 78, 14, 2, -23, 28, 16, -11, -3, 11, 66, 0, -20, 36, -16, -46, 32, 31, 29, 28, -45, -38, -4, -14, -49, 14, 6, 0, -63, -61, 5, 9, -16, 9, 57, -36, 7, -8, 28, -34, -16, -42, 10, -42, 12, -40, -26, -56, 29, -2, 10, 15, -2, -28, -21, -22, 39, 36, 59, -35, 27, 25, -16, -5, -32, 37, 15, -21, 10, -27, -23, 10, 40, -42, -38, 19, 38, 22, -15, 22, 45, -33, -19, -24, 34, -6, 46, -2, -21, 13, 25, 46, -15, 12, 22, 14, -34, 1, 55, -7, 46, -14, 1, -15, 29, -44, 19, -33, 26, 36, -4, -21, 14, 14, -13, -3, -32, 21, 0),
    (4, 13, -1, 9, -32, -34, -25, -14, -15, -10, -3, -28, 23, 21, 10, -41, -33, 25, 26, 14, 5, 18, 22, -23, 33, 3, 11, 51, 45, -7, 28, 29, 5, 18, 47, 36, 2, -5, 21, 6, 29, 50, -14, 5, 75, 15, -38, -10, 25, -24, -5, -10, 24, -11, 39, 7, 16, 18, 4, -11, -1, 3, -47, -28, 7, 5, -26, 10, 14, 4, 0, 4, 5, 16, -18, 3, -11, -43, 7, -1, 1, -24, -15, 16, 33, 89, 42, -1, 19, 26, -9, 11, 31, -17, 38, -48, 21, 18, -19, -1, 56, -9, 33, 37, -14, 24, 1, -15, 21, 82, -12, -28, 37, 36, 17, 22, 57, 39, 7, -46, 19, 44, 33, 17, 63, -41, 30, 25, -28, 11, 20, -16, 14, -2, 0, -5, 0, -36, -62, 16, 22, -9, -70, -4, -9, -45, -20, 27, -31, -28, -30, 5, -15, -17, 24, -22, 13, -15, 31, 35, 18, 0, 35, 1, 54, 9, 24, -12, -22, -8, -29, -1, 49, 6, 34, 17, -8, 53, 6, -4, -1, 48, 9, 39, 16, 21, -53, 49, -1, -14, -11, -13, -54, 23, 15, -38, 11, 7, 8, -29, -5, 17, -15, -18, 18, 18, -28, -16, -21, -7, -43, 28, -46, -36, -15, -7, -3),
    (3, 42, 17, 19, 31, -16, 6, 64, -49, -26, 0, -10, -18, 27, -14, 8, -11, -11, 4, 34, -9, -1, 1, 38, 3, 25, 16, 27, 60, -36, 32, 14, -19, 21, 1, -35, -3, 10, 8, 14, -17, 20, 2, -2, 7, 4, -22, -9, -45, -24, -18, -5, 35, 35, 34, 1, -35, 34, -31, -28, -38, -38, -45, -12, 8, -47, 4, 33, -9, -41, -20, -15, 27, 53, 0, 3, 21, 8, 25, 34, -28, -28, 28, 30, -50, 25, 19, -14, -33, -16, -21, 34, -22, -8, -14, 38, 19, -3, 64, 21, 51, -55, 52, 57, -37, 28, -34, 4, -69, -21, 20, -22, 10, -5, 27, 46, -7, 32, 14, 38, -6, -1, 5, -3, 2, -52, 2, -47, -22, 42, 18, 39, -14, -65, -46, 18, -37, -47, -25, -7, -10, -26, 16, -12, -18, -28, -39, 10, 34, -35, -24, 44, 10, -9, 25, -23, -42, 31, 1, 18, 7, 3, 20, -18, 46, 8, 7, -25, 31, 16, 5, 16, 51, 4, 39, 14, -54, 43, 13, 6, -1, 8, -34, 29, -49, -25, -21, 24, -4, 32, 50, 56, 34, -55, 23, -48, -3, -20, 22, -8, -16, 7, -15, 7, -42, -44, -4, 3, 8, -15, 24, -27, -23, -20, 30, 12, 2),
    (-40, -65, -27, 49, 21, -23, -51, -15, 7, -29, -50, 18, 35, 5, -53, 24, -4, -30, 15, 20, -3, -49, -40, -29, -32, -2, -20, 4, 49, -36, -97, -43, 30, -49, -27, -39, 16, -30, -27, -14, 7, -16, -11, 0, -20, -43, -29, -36, -18, 9, -18, -12, 9, -6, -79, -36, -44, -52, -8, -9, 16, -33, 37, 4, -9, -20, 29, -15, 6, -8, 18, -32, -51, 40, -19, 52, 13, -39, -29, -34, 31, 32, 19, -18, 58, -2, -19, -18, 16, 0, 39, 20, -3, -5, 7, -20, -41, -18, -34, 94, 8, -39, -44, 15, 25, -68, -45, 41, 73, -15, -29, -28, 11, -9, 21, 36, 50, 12, 9, -27, 30, -11, 13, 15, 4, 32, -29, -9, -42, -6, 28, 17, 8, 21, 46, 5, 30, 5, 43, 21, 58, -3, -19, 12, -29, 16, 28, -16, 17, 28, -8, 15, -37, 31, -15, -17, 8, 38, -7, -20, 8, -11, -40, -2, 0, -55, 50, 11, 48, 57, 20, -11, -9, -19, -21, 9, -7, -16, 27, -8, 6, 13, 28, -16, -31, -38, -16, 43, 5, 0, 30, 29, 31, 23, 20, 37, -13, 10, 13, 23, 25, 31, 14, -3, 45, 24, 9, -13, 23, -20, 5, 36, 40, 18, 23, 8, -6),
    (-29, 3, -30, 0, -14, -14, 0, 49, -51, 22, 0, 11, 31, -40, -32, -7, 37, -21, -6, 10, 21, 15, 29, 19, 2, -40, -3, 15, -61, -17, -13, 27, 17, -26, -22, 42, -16, -12, 26, 37, -11, -24, 5, -12, 32, -48, -12, -23, 30, 3, -14, 19, -8, 16, 30, 38, -18, 23, -48, 56, -2, 21, -33, 31, 44, 30, 55, -21, 38, -23, -5, -34, 44, -59, -25, 58, -16, -15, -9, 4, -54, -17, -37, 44, -18, 17, 25, 6, 7, -1, -15, -7, -40, -15, 6, 24, -17, -33, -52, 40, -3, 10, 3, -11, -30, -14, -45, 60, -14, -16, 27, -22, -14, -34, 6, -34, 28, -17, 17, -19, -2, -11, -38, 54, -15, -10, 9, 26, 12, 0, -48, 6, 63, -14, 41, 34, -21, 26, 46, -2, 31, -32, 20, -22, -16, -50, -61, -17, 40, 29, -9, -24, -60, -36, -3, -16, 7, 15, -34, 3, 7, -33, -7, -34, -32, 19, -35, -18, 9, -35, -62, 44, 62, -21, 6, -20, 0, -45, -21, -4, 14, -13, 6, -56, -33, -50, 16, 13, -7, -3, -16, -42, -16, 22, -29, 62, 28, 6, 5, -24, -15, -2, -67, 18, 47, -6, 8, -16, -17, -32, -14, 0, -21, -29, 41, -8, 2),
    (26, -52, -34, -5, -3, -11, -10, -9, -36, -11, -24, 32, 17, -28, -56, -34, 13, 4, -22, 18, -35, 8, -6, -1, 21, -3, 6, 18, 52, 5, 27, 7, 50, -6, 9, -49, -35, -77, -40, 10, 22, 30, 4, 5, -41, -31, -1, -26, -16, 26, 7, -48, -4, -12, 32, 45, 12, -48, 13, -15, -6, 27, -6, -66, 34, 23, -67, 2, -25, -27, -50, -8, -17, -3, 22, 29, 33, -32, 6, -28, -32, -46, -20, -24, 23, -11, 3, 33, 29, 33, 9, 21, -33, -14, 12, -26, -30, -16, 33, 58, -26, 15, 11, -17, 0, 0, -49, 18, 32, -23, -10, -16, -9, 3, 3, -48, 38, -2, -20, 35, -14, -1, 47, 27, 45, -9, 47, -63, -12, 44, -53, -9, 24, -14, -22, -40, 33, 2, -4, -17, 5, -32, 47, 25, -11, 18, -39, 14, 8, 36, -10, 3, 11, -29, -16, -29, 35, -32, -2, -8, 1, 23, -40, 9, -25, 26, -28, 38, 4, 14, -41, 12, -9, -23, 14, 11, -42, -18, -15, -15, -18, -2, -60, -58, 30, 16, -42, -41, -56, -21, 9, 58, 33, 24, 8, -23, 39, -20, 35, -23, -55, -20, -38, 35, -36, -46, -44, 15, -2, -32, 3, -12, -35, -34, 15, 44, -5),
    (-21, 23, -9, -34, 26, -17, 12, 1, 9, 38, -11, -30, -16, -20, 4, 2, -7, -5, -26, 12, 12, 40, -40, 57, -8, 27, -40, -43, -13, -18, -13, -7, -13, 30, 8, -13, 4, -29, -30, -21, 4, 19, -27, -50, -29, -51, -28, -8, -31, -34, -60, 42, -42, -39, 71, -39, -27, -57, -41, -8, -34, -1, 17, -44, -41, -13, 7, -73, -3, -8, 2, -2, -15, 41, 24, -33, 26, -39, 29, 19, 32, 38, 21, -44, 43, 17, -12, -6, 19, 29, -34, 31, 11, 15, -12, 48, -18, -7, -29, 9, 18, -44, -5, -26, -10, -6, -1, -40, 25, -13, -38, -43, -10, 29, 1, -39, -44, -55, 23, 99, -19, 43, 15, -4, 22, -13, 18, 7, -52, -37, -7, 45, -1, 3, 13, -37, 12, 19, 41, -61, -22, -49, 43, 45, -32, 19, 21, -50, 33, -46, -22, 1, -28, 24, 18, 6, -13, -20, -2, 5, -17, -44, -8, -7, -42, -30, -40, 24, -35, 8, -17, 0, 58, -15, -33, -4, -57, 24, 20, -9, -62, -34, 9, -12, 0, -9, 46, -14, -32, -13, -43, 3, 2, -22, 20, 9, 10, 32, -25, 16, -21, 10, -5, 31, 2, -7, 28, -39, 31, -17, 33, -19, 0, -55, 7, -3, -1),
    (-4, -32, -8, 46, 17, 0, 1, -17, -66, -40, -3, -34, -14, 3, 1, -32, 23, -34, -1, -63, 15, -23, -54, -4, 16, -33, -14, -16, 19, -39, 55, 19, -5, -57, 19, -21, 4, 18, -13, -33, 32, -39, -32, 18, 0, 43, 31, 40, -15, -5, -1, 23, 1, -27, 20, -3, -3, 22, 21, 12, -2, -4, 32, -34, 14, 29, 22, -44, -47, -22, 7, 47, -26, 25, -28, 45, 18, -44, 17, 2, -46, -35, 5, -29, -38, -36, -50, 1, 20, -19, 10, -27, -23, 26, 7, 14, 13, -10, 25, 24, -33, -44, 62, -23, -11, 13, -8, 27, -6, -29, -12, -55, -39, -34, 0, -5, -21, 47, -10, 52, 4, -7, 33, -18, 13, 39, 28, 40, -44, 29, 49, 33, 33, 2, 23, 7, 9, -41, 39, -9, -4, 35, 5, 18, 3, -59, -49, -41, 7, -7, 13, -47, -22, -1, 19, -27, -9, 43, -57, -28, 1, -32, -38, 6, -13, 37, 27, 39, 11, -29, 30, -11, 26, 24, 2, -32, -22, -12, -17, -5, -3, -4, -25, 1, -24, -11, 3, 24, -19, -2, 22, 4, -12, -15, 6, 32, -2, 30, 33, -6, -39, 27, 10, 6, 22, 43, -1, 10, 30, 6, 36, 9, -2, 17, 3, 22, -2)
  );
  ----------------
  CONSTANT Layer_6_Columns    : NATURAL := 8;
  CONSTANT Layer_6_Rows       : NATURAL := 8;
  CONSTANT Layer_6_Strides    : NATURAL := 1;
  CONSTANT Layer_6_Activation : Activation_T := relu;
  CONSTANT Layer_6_Padding    : Padding_T := same;
  CONSTANT Layer_6_Values     : NATURAL := 32;
  CONSTANT Layer_6_Filter_X   : NATURAL := 3;
  CONSTANT Layer_6_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_6_Filters    : NATURAL := 32;
  CONSTANT Layer_6_Inputs     : NATURAL := 289;
  CONSTANT Layer_6_Out_Offset : INTEGER := 3;
  CONSTANT Layer_6_Offset     : INTEGER := -1;
  CONSTANT Layer_6 : CNN_Weights_T(0 to Layer_6_Filters-1, 0 to Layer_6_Inputs-1) :=
  (
    (-4, -1, -16, 33, -7, -5, 33, 15, 0, -7, 29, -16, -20, 16, -4, -7, -26, 5, -36, 7, 5, 0, -31, -21, -15, -15, -31, 27, -37, -63, -10, -26, -15, -4, 28, 45, 4, -7, 37, 41, 22, -27, 24, -11, 28, 29, 39, 1, -28, 29, -27, -34, -1, 28, 12, 34, 28, -23, 16, 48, -9, -27, -7, -8, -36, -26, 21, 20, -22, -40, -29, 41, 27, -38, -41, -51, -32, 5, -37, -9, -4, -5, -31, -11, -28, 32, 22, 27, 50, 9, 7, 58, -51, -33, -17, 1, 14, 11, 31, 41, 3, 7, -18, 57, 5, 16, -26, -15, 41, -9, 48, 2, -13, 13, -43, -23, 4, 10, 19, 19, -24, 34, -19, 54, -23, 13, 21, -12, 44, 5, 34, 10, -13, 4, 3, 31, 1, 36, 30, -27, 42, -54, 40, 12, -14, 53, -41, -27, -24, -15, 34, -14, -9, 19, 10, -6, -30, 8, 0, -29, 19, 19, 29, 21, 8, -3, -14, 14, -20, 23, 22, -38, 44, -16, 26, 32, -17, 41, -20, -5, -10, -4, -8, -9, -24, -2, 13, 23, -12, -35, -26, -24, -22, 37, -1, -31, -36, -17, 24, 2, 25, -6, 0, 29, 36, -20, 9, -33, -9, 19, -1, 13, -21, 56, 30, -20, 3, 14, -10, 11, 37, 9, -40, -3, 1, 10, 27, -59, -43, -47, -3, 32, -40, -7, -31, 13, 25, -35, -16, -4, 2, -25, 1, 15, 13, 9, -15, -8, -19, -22, 6, 13, -17, 6, 3, 35, 50, 19, 21, -54, -12, -42, -53, 87, -51, 19, -39, -14, 16, -47, -40, 10, -19, -18, -8, -23, -38, -13, -43, -24, -45, -1, 1, -19, 3, -43, -8, -34, 2),
    (14, -13, 31, -19, 7, -18, -21, 24, -12, -11, 22, 27, 42, -37, -23, 44, 7, -17, 10, 16, -4, -5, -30, 0, -22, 17, 14, -6, -13, -18, -1, 30, 25, -5, -7, -6, 16, 8, -4, 4, 18, -3, -32, 12, 32, -55, -27, 35, -4, -13, 27, 30, 15, -4, -23, -27, -30, 14, 23, 20, -4, 2, -9, 5, -26, -2, 5, -11, 2, 5, 6, -58, -24, 23, -16, 2, 15, -34, 2, 32, 23, -1, 31, -25, 13, -17, 14, 11, 15, -27, 39, -19, -19, -29, -47, -4, 24, -36, 25, -15, 11, 8, 2, 26, -35, 32, -10, -24, -24, -17, -32, 57, 18, 18, -6, 36, 3, 7, -37, 19, -5, -22, 26, -1, -16, 11, 33, 35, -6, -17, 15, 8, -13, 37, -9, -50, -21, 26, -4, -4, -6, -36, -19, 52, 18, 11, -24, 38, -6, 34, -31, -29, 4, -14, 17, 18, -29, 33, -47, 21, 37, 0, 20, -51, -37, -2, 0, -72, -15, -13, 7, -5, -8, 7, -16, 47, -9, 9, 2, 25, 1, 62, -2, -34, -1, -43, 3, -23, -8, 37, 23, 5, 47, 0, 38, 19, 42, 38, 2, 41, 28, 7, 24, 1, 10, -59, -30, 14, -43, -5, -27, -18, 14, -34, -16, 12, -8, -27, 7, 17, -53, -13, -8, -14, 49, -24, 29, 22, 23, 12, -25, 14, -3, -2, 54, 26, -14, -40, -55, 9, 4, 17, -40, -3, 21, 19, 15, -25, -29, -36, 45, -5, -6, -21, 16, 5, 18, -6, -10, -25, -22, 31, -38, -8, 10, -27, 48, -1, -24, -1, -20, 32, 7, 19, -2, 4, -30, 28, -8, -13, 33, -16, 10, -13, -49, 33, -29, 41, -5),
    (20, 9, 26, -15, 2, 7, 0, 12, 31, -7, -8, -34, -12, 33, 1, -25, 41, -31, 25, -8, 44, -27, 15, -19, -21, -24, 14, -30, 19, 14, 14, -26, 12, 12, 26, 21, 1, 47, 8, 17, 16, 16, -11, -6, -14, 37, 33, -1, 42, 29, 14, -10, 21, -2, 35, 12, 22, 15, -2, -16, 24, 39, -2, -22, -28, 44, -12, 20, -7, 32, 4, -8, 35, -14, 19, 40, 12, 44, 59, 13, 43, 31, 9, -22, 15, 24, -26, -18, -3, 12, -14, 36, 37, 62, -20, 19, -18, -27, 52, 18, 6, 6, 11, -13, -27, 21, -19, 15, -24, 7, -40, 28, -11, 60, 2, 4, 17, 12, 9, -10, 13, -14, -15, 1, -21, 23, 53, 20, 20, 29, -17, -12, 20, 42, -32, -29, 4, -10, 10, 53, -26, -15, -13, 51, 10, 66, -37, 13, -16, 12, -16, -8, -12, -14, -31, -23, -2, 0, -5, 47, -10, 22, -15, -35, -27, 33, -8, -64, -4, -39, -5, 24, 15, 29, -24, 44, -5, 10, -5, 14, 15, -1, -26, -30, 25, -32, 26, -23, -26, -41, 6, 48, 18, -27, 51, -29, -8, 7, 12, 5, -22, 16, 15, 15, -2, 11, -34, 14, 0, 15, 18, -16, 14, -5, 24, 30, -39, -6, 19, 10, -23, -26, 4, 22, 0, 10, 23, -26, -20, -3, 4, -17, -33, -11, 8, 45, -22, 12, -7, -13, 6, 6, 18, -24, -15, 7, 11, -1, -8, 23, -6, -10, -34, -67, -15, 22, -13, 21, -5, -25, -19, -36, 1, -11, 9, 32, -5, 20, 18, 13, -13, -6, -29, -23, -2, 2, 7, -41, -13, -27, -30, 11, -12, -24, -30, -31, -31, 24, -5),
    (-26, -5, -16, 4, 0, -23, -26, -47, 24, -5, 45, 16, -5, -49, -13, 0, -1, -11, -11, 5, 9, -9, -21, -14, -3, 22, -5, -26, -15, -6, -32, -22, -26, 26, -14, -56, -19, -1, -19, 1, 0, -39, -20, -2, -13, -2, -44, 9, -12, 1, -3, -32, 28, 47, 32, 10, -10, -12, 27, -45, -4, 11, -26, -13, -1, -1, -36, -61, -27, -28, 1, 5, -20, 2, -7, -37, -27, -10, -55, 30, -62, 19, 8, -86, 3, 61, -8, -7, 14, 24, 26, -1, -14, -54, -48, -59, 0, -1, 2, -14, -57, 25, -40, 9, 7, 25, 8, 32, 14, -6, 11, -39, -9, -44, -19, -1, 13, -29, 11, 15, -11, -4, -42, 9, 38, -38, -60, -45, 18, 5, 36, -61, -8, -20, 5, 39, 27, 38, 5, -10, 6, -9, -10, -33, -9, 12, -31, -23, 4, -3, 29, 37, -5, 39, 13, -15, 1, -2, -25, 12, 49, 22, 30, -55, 35, -33, -20, 12, -24, 35, 32, -19, 44, -27, -65, -11, -45, -33, 8, -31, 0, -2, -48, 21, -8, -9, 57, 0, -18, -19, 8, 18, -32, -8, -16, 12, -20, 8, -70, -32, 51, -34, 7, -17, 4, 2, 23, 6, -3, 19, -10, -2, -25, -35, 6, -34, 13, -13, -39, -3, 26, -28, -77, -10, -4, 26, -9, 17, -6, 25, -46, -10, 3, 31, -38, 16, -4, -11, 6, -16, -16, 16, -32, 45, 36, -2, 21, 25, 27, -13, 5, 17, -6, -39, 2, -23, 3, 27, 36, -13, 56, 17, -22, 88, 30, 2, 8, 18, 26, -2, -3, 15, -39, 41, 7, -3, 27, -44, -22, 12, -40, 2, 3, -51, -20, -42, 18, 5, -3),
    (-41, -15, 21, -9, -33, -38, -16, -13, -3, 24, -21, -34, 14, 34, -31, -28, -38, -12, 9, -24, -25, 30, 1, -28, -11, -24, -30, -44, 32, -35, 13, -35, -54, 39, -28, -12, -17, -54, 34, 6, -30, -2, -66, -5, -23, -30, -63, -14, 9, -15, 18, -26, -26, -20, 13, 4, -18, -30, -52, -23, 7, -16, -15, 4, -19, 29, -14, 19, 19, 11, 26, -5, -22, -5, -35, 9, -19, 19, 17, -41, -2, 5, 27, -30, 9, -31, 21, -13, -25, -8, -22, 30, 36, 4, -2, 2, -72, 61, -3, -28, 7, -34, -2, -25, -31, -23, -36, -2, 46, 7, -25, -25, -30, -54, 33, -20, 8, 43, 0, -6, 3, -16, -36, -14, -18, -84, -24, -27, -51, 27, 15, -22, -9, -4, 20, 30, 5, 40, -14, -2, 30, -7, -25, -16, 2, -28, 42, 28, -6, -41, 29, 20, 2, 35, -10, 31, 0, -61, -18, -34, -31, -3, 23, -5, -6, 11, -12, 37, 17, 33, -4, 26, -2, 2, -18, -7, 24, -11, 4, 6, -12, 13, -20, 32, 9, 55, -18, 39, 25, -52, -11, -20, 1, 17, 7, 0, 21, -5, 50, 20, 3, 9, -41, -3, -11, -14, 24, -5, -7, -37, 43, 16, 14, 31, 23, 13, -25, 25, 39, 19, -1, -18, 15, 30, -1, 31, 30, -34, 29, -26, 41, 3, -17, 19, 21, 6, 33, -50, -24, -12, 16, -9, -21, -11, -10, 31, 4, 44, -18, -8, 24, 8, 14, 8, 33, -3, -11, -29, 17, -26, 25, 24, 13, 17, 27, -21, -19, 17, 5, 0, 36, 18, 25, 6, -5, 14, -1, 3, -15, 9, -20, 17, 16, 22, -13, 11, 1, 6, 0),
    (-45, 10, 7, -37, 8, 9, -19, -48, -19, -42, 31, -40, -7, -45, -16, 14, 23, 33, -29, -26, -30, 0, -12, -34, -5, -26, -24, -5, -7, 4, 18, 37, -42, -4, -26, 0, -13, 6, -32, -12, -26, -22, -33, -1, 18, 1, -27, 32, -21, -5, 2, -5, -24, 19, -3, -3, 24, -20, -21, -15, -35, -4, 38, 23, 8, 22, -42, 15, -26, 33, 46, 45, 2, -19, -44, -21, -9, 46, 5, -15, -14, -7, 25, 26, -17, 1, -34, 38, 4, -34, 6, 28, -42, 43, 24, 19, -42, -41, -38, -15, -28, -12, -32, 12, -21, -29, -40, -34, -32, -3, -32, -23, 0, -2, -19, 8, -12, 7, -53, 2, -17, -14, -25, 20, 10, -3, 30, -27, -20, 18, -41, -28, -11, -5, -8, -24, -2, -18, -70, -9, 21, -4, -19, 21, -3, -34, -26, -22, 9, 42, 1, -16, -29, 4, 31, 31, 3, -3, 34, -23, 23, -16, 8, -9, -6, -25, 43, -43, 4, -4, -54, -42, 35, -53, 27, 13, 24, -29, 2, 20, -32, 20, 26, 15, -14, -38, -7, 2, 19, -10, 8, 21, -2, 4, 22, 22, -41, -23, 20, 31, 0, -22, 28, -40, -34, 34, -16, 15, -20, 2, -37, -49, 14, 19, -33, -11, 34, 10, -22, 40, 25, -30, -4, 2, -16, 5, 30, -19, 33, -14, 10, 26, 18, -13, 6, 35, -33, 39, 13, 39, 30, -4, -15, 43, -11, 21, -48, 41, 35, 37, -3, 33, -12, 45, -1, 5, 0, -32, 32, -31, 21, 10, -5, -15, 29, -29, -18, 3, -3, -3, 45, 26, -16, -2, -29, 50, -11, 40, -5, 39, -16, -19, 6, -4, 30, 8, -29, -20, -1),
    (-35, 15, -9, 39, 12, -11, 15, 20, 37, 38, 0, -36, 26, 6, -9, -21, 39, -49, 32, 17, 0, -50, -7, 43, 10, -5, -29, 31, -12, 8, 20, -5, -22, -21, 30, -9, 8, -27, 2, 35, 26, -8, 7, -6, 20, 18, 22, -43, 40, -30, 24, 11, 7, -48, -18, 18, -46, 17, -16, 53, -4, 7, 15, -22, 29, -25, 15, -19, 39, -2, 62, -6, -12, 26, 1, 22, -9, -22, 19, -55, 15, 5, -25, -4, 4, -41, -21, 34, 16, -1, -9, -28, 2, -22, -11, 12, -2, -30, 25, 5, 13, -9, -2, -9, 21, 14, -21, -28, 14, -23, 11, -3, 12, 9, 53, 2, 11, 0, -5, 49, 10, 33, -40, 39, -20, 30, 63, 7, 8, -47, 42, 10, 21, 52, 44, 42, 34, -7, 26, -35, 30, -5, 9, 14, -25, 60, -20, -14, 43, 19, -9, 32, -9, 24, -20, 20, -1, 50, -16, 39, 26, 2, 7, 31, -10, 21, 37, 2, -15, -9, 1, -58, 6, 26, -11, -26, -13, 24, -40, -19, -15, 2, -8, 39, 27, -20, -4, -12, -79, 26, 4, -16, -50, 14, -6, 4, -33, 12, 6, -31, -16, 20, -32, -10, -16, -6, -31, -17, 17, 24, 25, 19, -26, -26, -26, -2, 9, -35, -23, 2, 16, -14, -17, 8, -26, 26, -34, -28, -37, -17, -17, -42, 17, 15, -13, -9, 36, 38, -16, 6, 18, 12, -10, 1, 17, 13, 16, -39, 11, -28, -26, 16, 14, -5, -16, -7, -41, -9, -30, -17, -19, -15, 32, -32, 18, -39, -22, 20, 37, 10, -23, 0, -22, -10, -24, 23, 0, 13, -22, 16, -7, -22, -5, 11, 18, 20, 51, -33, -3),
    (20, -17, -19, -23, -13, -35, 17, 6, -9, 6, 0, -56, 11, 2, -29, 28, -29, -4, 30, -6, -22, 31, -37, 32, -11, -11, -13, -57, 25, -31, 6, 34, 1, -4, 7, 20, -24, 10, -19, -21, -4, 7, 15, -25, -28, -18, -69, -3, -13, 46, 49, 10, -37, -46, 24, 19, -11, -53, -12, -37, 13, -19, 32, 37, -24, 21, -36, 54, 9, -14, 17, 6, 22, -44, 11, 24, 19, 30, -3, -10, -25, 2, 4, -14, -25, 12, -1, 14, -30, 0, -4, 23, -10, 7, -2, 28, 13, -16, -39, 11, 45, 26, 8, -1, -33, 24, 21, 25, -22, -16, -11, -23, -35, -38, 40, -40, -19, 1, -16, -5, -14, -42, 35, -14, -12, -49, 26, 8, -15, 23, 17, -33, -25, 11, 36, 2, -15, 0, 20, 11, 11, 0, -38, -8, -20, -27, 25, -36, -20, -39, -15, -35, -29, 30, 16, 21, 8, -48, 19, -19, -38, -37, -17, 10, 3, 11, -18, 41, 23, 22, -4, 8, 17, 12, 33, 6, -17, -53, 10, -3, 20, 28, -8, 11, -18, 41, -41, -19, 28, -58, -5, 11, -27, 0, -10, -11, -11, 10, 33, -1, 19, -8, 4, 24, -6, -48, -37, -6, -3, 16, 17, -31, -4, 27, 10, -6, -34, 5, -31, 28, 2, -37, 7, -35, 29, -18, -32, 13, -14, 26, -35, 23, 7, 26, 35, 23, 1, -11, -4, -30, -1, -11, -26, -13, 20, -10, 14, 58, -4, 22, 4, 18, -45, -8, -30, -22, 26, -33, 11, -13, 15, 37, 37, -16, 15, 24, 25, -19, 11, -28, 10, -11, -6, 2, 4, -30, -11, -32, -11, 60, 39, 10, 9, 38, -26, -5, 2, 26, 19),
    (-16, 27, -29, -22, 18, 18, 32, -4, -27, 21, -17, 6, -45, 7, -60, -13, -22, 3, 19, -18, -14, -44, 18, 42, 27, 39, -31, 24, 19, -21, 35, -10, -21, -21, 14, -11, 15, 17, 34, 22, 22, 2, 9, 22, 16, -36, -7, 17, -22, 7, 8, 12, 22, -34, -16, 33, -47, 33, 7, 17, 25, 14, 41, 24, 36, 20, -6, -36, -1, 14, 51, 7, 22, 0, -32, 15, 4, -8, 36, -6, 13, -10, 3, -8, 10, 19, -16, 12, -19, -8, 2, -20, 24, 7, 21, -3, 17, 30, 21, -37, 24, 33, 20, 14, -13, 10, 11, 5, -30, 2, -35, 37, -25, -25, -40, 15, 25, -55, 0, 58, 9, 33, -41, 32, -12, -11, 38, 40, 1, 7, 7, -31, 32, 8, -3, -15, 32, 0, 7, -1, 5, 30, -18, 29, 41, -10, -47, 17, 26, -35, 7, 44, -5, 39, 13, 60, -38, 24, 11, 18, 4, -50, -20, -17, 4, 14, 41, 19, -8, 20, 0, -13, 22, -22, 3, -37, -12, -6, -36, -4, -15, 8, 6, 19, -26, -9, 33, 10, -46, 19, 16, -34, -5, 19, -3, 15, 6, 16, -26, -33, 23, 3, 5, -14, 11, 41, -12, 25, -11, -11, -1, 13, -20, -15, -1, 37, -29, 25, 6, 43, -16, -49, 25, 25, -10, -12, 8, -14, -25, 16, 12, -9, -5, -35, -26, -14, -16, 57, 14, -24, 28, -5, 13, 17, 16, -10, 10, 51, 28, 6, -28, 6, -9, -6, 29, 29, -48, -25, 15, 40, -2, -18, -3, 3, 16, -24, -1, -48, 17, 9, -13, -19, -27, 7, 7, -9, -19, 27, 22, 44, -12, 17, -20, 35, -56, 15, -20, 25, -6),
    (5, 36, 15, -48, -5, -5, -8, -72, -24, 3, -12, -34, -26, -55, -32, -22, -33, 8, -92, 38, -32, 20, 6, 24, -35, -10, -18, 9, -29, -44, -24, 27, 17, 9, -8, -2, -4, -29, -17, -10, -21, -14, -44, -23, 1, -14, -12, 25, 33, -15, -36, 26, -33, 1, 34, -20, -23, 7, -13, -11, 2, -1, 39, -5, -8, -10, -34, -6, -29, -31, 4, -41, -6, -9, -48, -44, 2, -7, -27, 21, 30, 39, 9, 24, -23, 1, 22, -3, 0, -38, -16, 34, -1, 1, 4, -2, 41, -4, -5, -16, -16, -18, 42, 43, -18, -12, 21, 43, -6, -10, 49, -8, -17, -13, -35, 22, 7, 50, 5, -20, 11, -1, -4, -5, 9, 7, -12, -12, 33, -18, 44, -23, -28, -7, 37, 0, 33, 18, 12, 22, -20, 5, 33, -13, -20, 1, -53, 20, 37, -8, 35, -6, -17, -15, 6, 1, 26, 17, 21, 25, 48, 8, 28, -23, -6, 21, 23, -16, 13, 31, 28, 3, -47, -19, 11, 45, 2, 20, -34, -19, -9, -18, 25, -22, 5, 11, 57, -14, 5, 18, -53, 26, 30, -26, 2, -7, -22, 45, -22, 33, -9, -39, -12, 19, 8, 17, 36, 5, -11, -42, 2, -39, 0, -37, 0, 5, 16, 7, -21, -26, 3, 0, -5, 25, 28, -5, 16, -14, -30, 41, -13, 14, 30, 5, 48, -21, -10, 2, -1, 26, -39, 32, -16, 4, -22, -44, 17, -6, 17, -6, 23, -33, -12, 32, 14, 20, 34, 5, -2, 8, -3, 19, -13, -8, 7, -17, -5, 25, -16, 44, -15, 18, -23, 9, -35, 8, -37, 7, 3, 8, 25, -3, -2, -11, 20, 37, -11, 4, -5),
    (1, 26, -58, 1, -46, -52, -22, -45, -5, -6, 8, 26, -1, 18, -12, 14, -14, -46, 11, 21, 6, 2, -30, -3, -2, -17, 26, -54, 41, -44, -11, 10, 4, 26, -41, 5, -17, 10, -32, -23, -10, -10, -29, -14, -12, 36, 19, 0, -1, -31, 28, 7, -20, 8, -9, -16, 26, 28, 2, -20, -17, -9, -14, -65, 37, -38, -20, 18, 47, -41, -30, 24, -5, 2, -41, -55, 50, -20, -1, 1, 8, -31, 4, -5, 28, 5, -1, 42, -4, 15, 62, 16, 18, -11, -17, 1, -25, -35, -52, -29, 11, 11, -6, -8, -10, -12, -24, -12, 35, -2, -29, -27, 21, -19, 66, -24, -48, -10, 19, 13, 0, -4, -15, -12, 8, 15, -12, -39, 46, -43, -1, -12, 45, -21, 12, -4, -10, 10, 1, 24, -3, 8, -6, -11, -7, 17, 43, 1, -17, 25, 23, -11, -31, 40, -11, -37, -27, 3, 15, 26, 17, -12, 25, 5, 59, 19, -1, 15, 41, 3, -13, -43, 8, -5, -5, -25, 16, -5, 22, -17, 2, 26, -19, -25, 0, -31, -11, 7, 13, 19, 24, 3, 50, 22, 10, 0, 39, 28, -12, 23, -21, -19, 12, 19, -1, 5, -18, -31, 3, 1, 7, -25, 12, -21, 33, 0, 15, 18, -16, -14, -16, 13, 7, -22, 14, -6, 37, -9, -1, 20, 21, 34, 11, 35, -11, 25, 24, -40, -5, -35, -4, -4, 38, -33, -23, -45, -30, 42, -29, -24, 12, -31, -22, -33, 32, 8, -52, -11, -34, -36, -3, -12, 16, -4, -32, 36, 11, -30, 6, -3, -18, -51, -6, -61, 7, -56, -31, -1, 3, -20, -10, 0, 12, -38, 22, -3, 23, 9, 16),
    (-1, -43, 17, 14, 38, 21, 52, 24, 10, 35, -7, 14, 25, 12, -17, -8, 4, 7, -65, 11, 6, 43, -15, -12, 40, 7, -8, 57, -22, 18, 0, -20, 27, -37, 36, 30, 21, 19, 58, 60, -7, -9, 34, 20, 39, -3, 27, -3, 11, 11, -27, 23, 31, 28, -2, 29, -10, 16, -8, 38, -27, 28, 10, 15, -9, -45, 20, 7, 39, -5, 57, 5, 17, 38, 34, 8, 5, 31, -30, 0, 0, -3, 21, -18, 26, 44, 8, 0, -34, 16, -20, 34, -24, -7, -37, 35, -23, 1, -5, -25, -35, -10, -30, -35, -21, -53, -38, 31, 14, 27, -22, -23, -47, -7, 20, 8, -40, -32, -41, -12, 21, 10, -55, -9, 14, -8, 55, 50, 17, -35, -12, 51, -41, 36, -24, -38, 34, 30, -18, -30, 48, -1, 17, -16, -19, -10, 44, -1, 12, -22, 0, -15, 26, -18, -39, -29, -39, 19, 33, -4, 30, -3, 22, 25, -19, 30, 4, 41, 13, 11, 6, -33, 40, -18, 13, 28, -36, 2, 24, -32, 32, 2, 15, 5, 33, 9, 14, -8, -27, -3, 10, -8, -16, 10, -12, -45, -21, -20, -18, -49, 5, 18, -2, 3, -7, 14, 25, -15, 8, -58, -3, 24, -42, 15, -29, -32, -4, 3, 7, 30, -1, -39, -1, -15, -33, 47, 18, 2, -25, -16, 21, -21, 2, -25, -28, -3, -41, -53, -15, 9, 10, -51, -21, 9, -33, -34, -5, -13, -23, -26, -2, 5, -8, -12, 4, 7, 13, -7, -34, 7, -18, 24, -47, -27, -33, -20, -20, 24, 28, -26, -23, 27, -17, -54, -21, 2, -25, -32, 25, -20, 19, 34, 5, -11, -3, 8, -39, 25, 5),
    (-7, 27, -16, 18, 37, 11, -43, 52, 26, 22, -37, 14, 24, 10, 2, -18, -21, -38, 19, 6, 18, -23, -19, -4, 18, 3, 10, 51, 21, -4, -17, 31, 23, 0, -11, -12, 24, -29, 10, 24, -13, -10, 2, -23, 16, -37, -22, 22, 4, 26, -32, 29, -33, 12, -11, 30, -49, -7, -10, -20, -21, 14, 39, 33, -17, 29, -39, -33, 15, -18, 14, -4, -35, -18, -42, -23, -24, -66, -24, 20, -5, 15, -1, 24, -43, 7, -9, -24, -35, -26, 6, -28, -26, -29, 43, 39, -25, -47, -15, -23, 3, -25, 36, 36, -9, 13, -40, 32, 24, -8, 6, -28, -27, -46, 5, 16, -30, -8, 3, -35, 14, -15, -24, -22, -24, -27, 32, 28, -16, -14, -28, 30, 19, -35, 83, -1, 15, 46, -31, -2, 15, 22, -30, 30, -21, 6, -27, -14, -8, -8, -38, 15, 14, -21, 24, 11, 45, 38, 37, 23, 2, 35, -10, 35, 20, 31, 62, 34, -42, -18, -62, -22, -40, 21, -29, 19, -35, -42, 30, 22, -12, -21, -15, 18, 24, -34, 36, 9, 39, -9, 32, 17, -14, -30, -12, 19, -50, -2, 23, 18, -3, 2, 17, -41, -5, -33, 35, 20, -24, -41, 5, 18, -39, -9, -15, -25, 25, -20, 5, -42, -47, 8, 19, 18, -5, -7, -21, -22, -60, 30, 49, 43, 36, -6, 14, -27, 21, 0, -27, -19, -36, 10, 46, -48, 27, -25, 11, 14, 15, 42, -18, 7, 27, 20, 6, -24, 22, 19, 24, 38, 19, 30, 34, 49, 41, 40, 6, -13, 1, -24, 6, 2, -6, 16, 46, -46, 18, -10, 5, 17, 1, -13, 6, 13, 34, -14, 23, 13, 5),
    (-23, 15, -3, -29, 28, -3, 9, 12, 18, -26, -24, -7, 1, 31, 40, 7, 32, -19, -38, 43, 42, 8, 28, -2, 20, -3, -9, 54, 32, 21, 4, 37, 21, -29, 35, -19, -37, 37, -21, 20, 15, 3, -19, 0, 35, 1, 29, 39, 40, 19, 11, 0, 48, -5, 39, 11, -28, -18, 18, 44, -5, 41, 29, 22, 49, 4, 15, 10, -23, -10, 7, 42, 22, -28, -6, 31, -16, -37, -4, -15, 15, 12, -16, 14, -3, -29, 5, -16, -60, -10, 20, -44, 24, 16, 40, 43, -16, -44, -51, 25, -31, 1, 16, 0, 7, -2, -28, 3, 4, 41, -4, 4, -3, -10, 11, 9, -30, -5, -41, -31, 12, 20, -35, 9, 16, 32, 40, 12, -4, -41, -9, -15, -32, 50, -4, 12, -6, -13, -35, 18, -11, -27, 37, -19, -6, 17, -14, 8, 8, -5, -22, -26, 12, 20, -24, -48, 13, 54, 23, -17, -11, 9, -24, 47, 0, -22, 25, 25, -6, -16, 20, -11, 2, -52, 22, -33, -4, 13, -32, -48, -32, -27, 8, -1, -11, -18, -19, -44, -33, 6, 22, -24, 13, -63, -27, 33, 6, 40, -24, -3, -29, -37, -7, -2, 30, 30, 4, -29, -11, -16, -70, 16, 4, -20, -22, -32, 54, -28, -36, 42, -12, 28, 30, 13, -13, -44, -14, 40, 13, 2, -12, -31, -2, -29, 8, -3, 20, 26, -24, 23, -22, -3, -12, -21, -3, 40, -17, 14, 7, 16, 24, 30, -24, -21, -33, 9, 23, -40, -8, -22, -3, -17, 16, 16, 20, -18, 45, -22, 27, -6, -47, 9, -26, 9, -23, 5, -4, 6, -20, 43, -34, -8, 48, 17, -41, -12, -1, -27, -19),
    (17, 28, 8, -9, -32, 51, -41, -59, -25, -7, 23, 10, -1, 6, -10, 3, 24, 27, -7, 2, 14, -7, -34, -54, 1, -29, 27, -28, 21, 2, -28, 54, -15, 46, -23, 45, -52, 5, -35, -35, -2, 6, -5, 5, 23, 30, 28, 27, -37, -3, 28, -4, -26, -17, -6, -13, -22, 6, 41, 17, -18, -4, 21, 37, 7, 5, -20, 34, -7, 9, 16, 15, 7, -12, 8, 7, 36, -57, 44, 45, 5, -61, -28, -70, -41, -23, -57, 9, -11, -15, 18, -26, -37, -14, -24, -20, -24, 23, 14, 11, 7, 23, -35, -1, -55, 0, -14, -14, -4, 2, -27, 22, -3, 9, -55, 28, -26, 21, -19, 14, -50, 16, 15, -13, 20, -21, -20, 37, -35, 28, -57, 21, 16, -53, 4, 10, -23, -26, -4, -13, 2, -1, -34, 6, -23, -27, 28, 27, 14, -13, -8, 20, -35, 16, -7, -30, 11, 1, -4, -46, -28, -30, -1, 14, 13, -25, 30, 10, -26, -9, -14, -54, 2, -6, 23, -4, -33, -13, 25, -5, -36, 1, 14, 26, -14, 5, -8, 3, -10, 29, 18, 15, -9, -27, 36, -20, 3, 5, 14, 36, -50, -6, 7, 22, -12, -6, -10, 46, 4, -19, -10, 24, -33, -1, -6, -12, -5, -15, 11, 32, -40, 39, -36, 28, 3, 44, -17, 8, 12, -37, 12, 12, 16, 7, 4, 41, -26, 49, -55, -7, -13, -15, 1, -6, -20, 30, 28, 29, 17, -16, -10, 19, 12, 23, 22, -12, -34, 7, 31, 16, 26, -18, 0, -6, 10, 29, 0, -29, -2, 25, -30, -60, -13, 8, 28, 31, -9, -28, -9, 14, 4, -19, 0, -1, -22, 23, 33, -3, 27),
    (-16, 28, -41, -59, 5, -42, -1, -44, 30, -7, -29, 19, 2, -16, -30, -37, 23, -30, -37, 12, 6, 22, 29, 10, 34, -10, -34, -17, -23, -24, -36, -1, 5, -28, 23, -2, -27, -12, -20, -10, -4, 34, 19, 9, 4, 26, 0, -7, -1, -21, -8, -21, -20, -37, 8, -13, -2, 41, -32, 42, 11, 15, -3, 29, -53, -31, 20, 32, -58, -33, -5, -20, 26, 13, -48, 1, -6, -33, 15, -54, 3, -43, -33, -26, 41, -27, -38, 36, -20, 26, -7, 7, -11, -15, 12, 22, -22, -12, 15, -44, 21, 31, -1, -1, -60, -15, -35, -11, -45, -26, -23, -19, -29, -48, -32, -34, -36, -56, -56, 6, -23, -38, 16, 23, -44, -9, -19, 28, 31, 22, -5, -22, -6, 41, 23, -25, -15, 43, -3, -30, 24, 2, -32, -1, -6, 29, -33, 14, 37, -62, -10, -4, 4, 24, -13, -21, -34, 7, 1, 14, 14, 28, 5, -5, -4, -10, -18, -3, 46, -11, -33, 13, 26, 18, -37, -8, -9, 20, -33, 28, 38, -52, 24, 26, -35, -6, 11, 45, -3, -22, 10, 20, -30, 11, 6, -7, 21, -6, 51, 18, 0, 22, -20, 13, 23, 14, -2, -37, -37, -26, 11, -8, -7, -12, -36, -6, -17, -20, -7, 49, 38, -11, -13, -21, 20, -13, 3, -24, -10, 37, -6, 21, 24, 37, -4, 5, 10, -42, 39, 18, 0, 0, -2, 22, 13, -8, -15, -10, -39, -5, -24, 2, 12, -21, -21, 42, 9, 14, 22, 4, -19, -19, 3, -3, 33, 27, -6, -11, 29, 10, 26, 25, 25, 13, -32, -3, -16, -49, 37, 19, -21, 2, 14, 17, 1, -7, 13, 48, -3),
    (13, 9, -36, -31, 7, 40, 13, -32, -23, -12, 8, 51, -45, 16, -32, 16, -25, 0, 19, 7, -32, -3, -16, 4, -16, 5, -11, -57, 12, 19, 17, -14, 19, -10, -5, -19, 16, 32, -27, -2, 18, -13, 47, 52, -10, -22, 11, 39, -15, 14, -10, -28, 1, -39, -32, -45, 0, 12, 16, -64, -33, 21, -33, 27, 19, 33, 2, -45, 10, 33, -51, -9, -21, -19, 43, 42, 0, -44, 34, 31, 42, 22, -26, -33, -1, -54, -3, 5, 36, 8, 21, -54, 37, 24, -27, 43, 16, -16, -36, -25, -4, -18, -35, -12, 12, -21, 39, 42, 33, 27, -17, 18, 12, -14, 44, -1, 23, 39, 8, -22, -3, 47, 17, 29, 16, -42, -10, -38, -16, -27, -26, 2, 11, -9, 26, -18, 5, -18, 39, -3, 35, 5, -28, 8, -23, -20, -26, -5, 25, 6, -8, 33, 21, 43, 13, -13, -21, -63, -2, -25, 1, -23, -15, 41, 16, -1, -23, -15, -8, -14, 40, -28, -26, 6, -18, 53, -4, 19, -15, -1, -10, -31, -62, -26, -25, -1, 36, 0, -17, -45, -25, -25, -1, 28, 0, 13, 39, -32, 0, -30, -2, 15, -12, 35, 8, 6, 35, 40, 6, 42, 6, -19, -17, 40, -53, -23, -13, -5, 29, 38, -20, -13, 11, -37, -23, -59, -25, -25, 20, 6, 6, -53, 18, -23, 19, 17, -12, 8, 26, -43, -29, -17, 9, 7, 15, 34, -25, -10, -1, -19, 32, 23, 10, -6, -35, -6, -6, -5, 6, 36, 19, 46, -15, -22, 16, 7, 60, -10, 5, 31, 14, 18, 12, -23, -33, 7, -35, 20, -2, 10, 7, -45, 12, 32, -25, -34, 1, -4, 5),
    (-31, -19, 39, -23, -54, -41, 34, -39, -21, -37, -46, 6, -9, -30, -44, 61, -60, 33, -25, 45, -15, 49, -14, 9, -43, -1, 37, 20, 24, 54, 20, 25, -32, -1, -8, 1, -37, -7, -42, 6, -26, 36, 6, 3, -29, -51, -61, 18, -36, -27, 29, -28, -25, -44, 5, 0, -17, 40, 8, -12, 13, -47, -52, -24, 31, -10, -1, 23, 42, -17, -13, -18, -10, 48, 15, -21, -1, -45, -19, 12, 47, 8, -49, -15, 4, 9, -8, 29, -13, 49, 24, 26, 2, -17, -28, -52, -10, 34, 20, -44, -41, -18, 20, -35, -23, -10, -20, 22, 6, -41, -22, 19, 6, 23, 5, 31, 10, 44, -14, -6, -29, 3, 42, -8, 40, 57, -6, 4, -12, -17, -21, -15, -17, -48, 3, -6, -48, 30, -49, 22, 9, -1, -14, 44, -8, -16, 37, -8, 24, -33, -12, -14, -15, 32, 35, -13, 15, 34, 2, -44, 10, -22, -10, 30, 44, -10, -6, -4, -13, -6, 0, -7, 9, -72, -1, -10, -5, 39, -19, -44, -9, -15, 0, -12, -33, 6, 30, -26, -58, -3, 0, -21, 5, 12, 4, -26, 31, 1, 2, -28, -24, -1, -4, 26, 27, 13, -5, -27, 35, 40, -26, 14, 20, 19, -17, 38, 10, -20, -1, -9, -8, -6, 18, 1, 11, 34, 16, -23, 17, -35, 6, -56, -30, -20, -44, 2, -11, -15, -11, 19, 2, 39, -4, 50, 11, 44, -10, 20, 9, -28, -20, -3, -13, 4, 9, 13, -39, -24, 19, 4, -37, -22, 9, -46, 11, 33, 1, -32, -43, 33, 5, 7, 18, 21, -65, -12, -5, 31, 50, 14, 16, -46, 12, 20, -17, 56, 1, -1, 8),
    (-47, -37, 27, -20, 27, 24, 22, -27, -27, 6, -15, 2, -7, -42, -46, -17, 45, -4, -15, -18, -13, 5, -36, 27, 1, -10, -25, 57, -22, -5, -1, 4, 11, 10, 42, -7, 16, 26, 35, 8, -18, 18, 34, 5, -6, -55, 8, 12, 32, 23, -81, -6, 20, 6, 22, 23, -14, -6, -44, 46, 10, -22, -23, -3, 7, -9, 12, -53, -22, 10, 11, 20, 5, 47, 26, 11, -10, -36, 54, 4, 4, 1, -84, 17, -5, -30, -30, 21, 5, 9, 23, 17, -38, -5, -34, 23, 15, -53, 43, -2, 57, 4, 14, 21, 9, -9, 14, 15, 21, 24, 14, -25, -29, 6, 23, -18, 15, 33, -37, 39, 35, 29, -50, 32, -18, 51, -5, 20, 0, -2, 23, -30, 46, -4, 47, -36, -41, -22, 34, 2, -24, 10, -11, -19, -30, 66, 30, -16, 21, -29, -3, 32, 8, -11, 8, -11, -49, 41, -17, 14, 37, -23, -16, -43, -14, 10, 40, -6, -30, -39, 43, -6, -43, -4, -27, -7, -15, 29, -60, -7, -15, -38, -26, 13, 25, 9, -2, 0, -43, 7, -47, 35, -42, -41, -25, -29, -3, 7, -11, 27, -26, -35, -2, -12, -41, 16, -5, -26, 54, -51, -21, 0, 1, 13, -33, 16, 27, 1, -29, 25, 30, -11, 2, 16, 0, -30, 26, -36, 12, -43, 38, 4, 23, 6, 32, -14, -15, 33, 20, 1, 10, -54, 15, -40, -7, -9, -20, 4, 26, 0, -59, 46, 3, 18, 35, 8, 14, -29, 14, 21, 14, -30, 29, 34, 46, 10, 10, 17, 0, -12, 26, -45, -8, -34, -16, -27, -18, 47, 26, -25, 16, 9, -22, 38, -21, -4, 39, 5, -2),
    (10, -39, 0, 22, 77, 1, 9, -15, 16, -34, 8, -30, 60, -42, -42, -31, -17, -46, 50, -30, 27, 14, -15, 2, -40, -14, 1, -35, -47, 0, 2, -11, 13, 7, 5, 22, 32, -42, 30, 50, -29, -1, -59, -18, 22, 7, -30, 7, -44, 4, 10, 23, -18, -37, -4, 1, -7, -30, 23, 29, -33, 5, 56, 35, 7, 18, 13, 13, 4, 37, -22, -24, 16, -20, -18, -44, 34, 8, -52, -8, -37, 27, 2, 18, -28, 15, -29, 14, -37, 28, -27, 14, -25, -13, -8, 8, 25, 6, -35, -28, 16, -29, 81, -35, 5, -43, -25, -49, -15, -27, 16, 15, -22, -33, -20, 24, -33, 42, -31, -12, 17, -30, -24, -15, 32, 24, 45, -18, -36, 2, -10, -22, 3, 17, 23, 15, -37, -4, -38, 1, 19, 12, 5, 8, -30, 10, 50, -11, -48, 2, 22, 25, -16, 50, 16, 21, -16, 29, 25, 22, 2, -3, 24, -15, -14, 36, 35, 0, -17, -9, -34, 24, -31, 22, -54, 31, -23, -4, 4, 9, 7, -48, 1, -4, 0, 45, -8, 33, 18, -26, 33, -4, 5, -9, -19, -36, 1, 16, 47, 17, -12, -12, 1, 19, -45, -24, -13, 1, -10, 16, 51, -26, -23, -29, 21, -7, 15, -20, -26, 5, -6, 33, 54, 30, -16, 34, 16, -39, -21, -12, 8, 2, 8, 3, -19, 2, -5, -56, 40, 32, -42, 8, 28, 18, -5, -12, -14, -18, -35, 48, 3, 44, 35, -29, 49, 20, 1, -10, 22, -13, 7, -26, -22, 29, 21, 41, -32, -8, -18, 15, 0, 2, -12, -17, -10, 24, -23, -13, 22, -19, -38, 43, 13, -4, 26, 14, 14, -25, 4),
    (-11, 8, -33, 16, 8, 20, -3, 19, -9, -43, 12, 4, 20, 23, -13, 18, 17, 19, -53, 4, -27, 46, -19, -42, -13, 17, 26, 34, -4, -21, -44, -21, 0, -36, -3, 27, 42, -34, -40, -26, 20, -20, 5, -42, -22, 5, 8, -16, 5, 14, -32, -11, 8, 30, -28, -12, -15, -13, 10, 28, 10, -36, -11, -26, -1, -32, 24, -7, 38, 15, -16, 22, 18, 18, 6, -11, -2, 3, 10, 32, 27, 26, -17, -14, -11, 43, 0, 11, -9, -19, -23, 5, -41, 38, -19, -37, 10, -7, 6, 11, -12, -1, -5, -21, -35, -6, -19, 4, -7, 12, 21, -28, -11, 14, -32, -5, 40, 11, -8, -36, 20, -44, -8, 20, 30, -12, -43, -4, 16, 12, 45, -14, 10, 16, -49, -35, 27, -27, 20, 12, 25, -37, 12, 37, 40, 22, -9, 30, -10, 40, 43, -28, -22, -3, -10, -28, 8, -10, 2, -25, -24, -6, 27, -39, 12, 7, 6, -4, -16, -22, -22, 9, -13, 8, 18, 10, 1, 12, 7, 55, -2, 37, 37, -24, -28, 0, 7, 25, -8, 9, 21, -4, -58, -14, 8, -47, -14, 26, -6, -15, -43, -48, -11, 31, -67, 28, -17, -44, 14, 2, -7, 12, 9, 6, 19, -34, 0, -61, 7, -46, 23, 40, 9, -34, -29, 16, -5, -64, 1, 10, -57, -20, 17, 36, -40, 12, -2, -27, 29, -21, 25, 34, 27, 20, 9, 13, 14, -47, 8, -28, 7, -58, 28, -24, -15, -28, -13, 16, 32, 34, 37, -3, -4, 24, 2, -14, -55, 9, -19, -24, 16, -14, 39, -4, -34, 10, 12, -29, 30, -22, 2, -1, 4, -5, 14, 27, 39, 27, -7),
    (33, 15, -33, 26, -25, -27, 2, 14, 24, -31, 6, -18, 21, 57, 19, -4, 11, -22, 35, -44, -6, 26, 25, -15, 36, -31, -54, 2, 4, 40, 17, 9, -41, 15, -8, 34, -18, 12, -13, -22, 34, -45, 28, -14, -11, 4, 8, -1, -9, 19, 23, 15, -13, 49, 7, -45, -7, -18, -53, -20, 19, 34, -11, -21, -34, -34, -8, -13, -17, -23, -16, -25, -14, -35, -19, 32, -6, -16, 5, -22, 14, 6, 20, -4, -5, -9, -17, 6, 15, -6, -6, -10, -11, 4, 11, 25, 2, 15, 21, 61, -35, -6, -9, -41, 58, -38, 11, -45, 21, 20, 58, -23, 46, 31, -1, -4, -2, -12, 17, 30, 26, -8, -23, 5, 10, 15, 17, -19, -11, -5, -3, 18, -34, 18, -26, 2, 19, -5, 26, -55, 6, 40, 48, -9, 15, 44, -22, 29, -21, 17, 27, -8, 57, -14, -31, 46, 0, -6, -20, 20, -21, -41, -40, -37, -53, -35, -6, -49, 16, -41, -30, 34, -22, 8, -39, 11, 2, -21, 21, -15, -46, -13, 3, 20, -6, -30, -27, -39, -27, 6, 10, -22, -12, 11, 4, -18, -22, -27, -5, -6, -3, 27, 21, -21, 21, 48, -28, 6, 36, 35, -22, 27, -18, 0, 43, 30, 3, -21, -3, -31, 29, 8, 10, 17, -8, -6, 33, 51, -16, -24, -24, -34, -1, 19, -20, -15, -26, 10, -4, -9, -2, 20, -2, 47, -9, 0, 7, 32, 52, 4, -47, 15, 21, -19, 0, -6, -36, 26, 20, 20, -30, 1, -14, -5, -18, -3, -31, -3, -27, 53, -40, -26, -28, -26, 32, 20, -30, -11, 1, 30, 34, 19, -14, 3, -4, -27, 9, 15, -1),
    (-18, -32, 8, 4, 24, -29, 20, -17, 26, -23, 8, -15, 34, -30, -36, 19, -9, 7, -2, -50, -17, 44, 17, -24, -9, 29, 0, 20, -1, -28, -41, 30, -10, -32, -3, 31, 25, -41, -26, -16, 16, -7, 5, -17, 28, -1, -40, 11, 6, -9, -29, 2, -32, 53, 16, -6, 11, -35, -35, 44, 33, -19, -27, -9, -44, 9, 16, -38, -15, -20, -1, -41, -6, -2, 9, 6, -16, 30, -56, -22, -15, -26, 9, 41, -16, -4, -5, 14, 24, 4, -21, 15, 10, -45, -30, 7, 35, 2, 24, 69, 35, 31, -20, -12, -24, -13, 43, 37, 33, -2, 22, 7, -1, -19, -17, -3, 22, 25, -23, -38, 19, -12, -3, -43, 24, -10, -40, 28, -17, 13, 20, -16, -4, -2, 21, 30, 17, -14, 14, 15, -1, -12, 36, 5, -24, -7, 4, -10, 25, 9, -10, 14, 10, 13, 1, -24, 9, 10, -2, -2, -2, 44, 36, 7, -26, 23, 26, -1, -10, -17, -17, -15, -2, -10, 31, 39, -28, 14, 6, 7, 17, -9, 3, 7, -40, 0, 42, 18, 5, 8, -35, 9, -32, 6, -39, -5, -47, -54, 8, -2, 39, -8, -26, -5, 16, -10, 17, -21, -15, -35, 24, 7, -28, -9, 44, -8, -14, -5, -43, -28, 0, -28, -27, -12, -49, 48, -39, -67, -26, -12, -20, 23, -13, -15, -72, 13, -7, -4, -33, 6, 15, -12, 62, 12, -37, -14, -16, -9, 17, -11, -16, 1, 12, 2, -15, -39, 37, 45, 5, 28, 29, -27, 21, 53, -32, 30, -62, -23, 45, -40, -21, 40, -5, -25, 14, 5, -11, -16, -28, 16, 42, -19, 41, 11, 32, 28, 54, -7, 11),
    (0, 13, 23, -3, -39, -15, -21, -3, 0, -21, 15, 27, -40, -15, -21, -14, 12, 33, -86, -18, -4, -25, -8, -19, -18, -17, 0, -2, -6, -17, -52, 0, -1, -19, 15, -20, 24, -33, -52, -23, 21, 20, -41, -2, 41, -5, -22, 20, -30, -27, -7, 13, 2, 10, -31, 25, 31, 26, 33, -16, -32, 27, 18, 22, -15, -58, -12, -8, 41, 16, 55, -16, -18, -23, -46, -56, 55, 5, 10, -42, -22, -51, 11, -39, -42, 8, -26, 38, 33, 20, -5, 24, 4, -16, 9, -20, -1, 14, -29, -3, -61, 15, -11, -3, 16, 9, 21, 19, -33, -19, -25, 4, 29, 28, -43, -15, 4, -17, 19, 11, -3, -6, -38, -22, -32, 7, 12, 35, -1, 3, 22, 10, 23, -15, 16, 34, 18, 37, -16, -2, 37, -47, 5, 6, 28, -30, -25, 36, -49, -76, -27, 24, -33, 27, 8, -8, 37, -34, 39, 15, -9, -8, 2, -1, 37, -45, 2, -12, -2, 22, -63, -15, 26, -3, 17, -38, 10, -23, 34, -21, -16, -41, -11, 56, 0, 26, 6, -7, -19, -24, 70, -13, -10, -26, 0, -15, 10, -21, -66, 39, 35, -2, 26, 14, 41, -44, 11, 19, 41, -29, -14, 22, -10, -38, -5, -4, -52, 44, 4, -3, -9, -28, 11, -6, 3, -13, -6, -11, -13, 16, -36, 29, 6, 5, -43, 41, 3, -22, 4, 15, 26, -4, -6, 2, -6, -12, 13, 19, -36, -17, 4, 26, -9, 16, 9, 21, 1, -18, 19, 6, -7, 14, -17, 22, 17, -5, -28, 1, 34, -5, 23, 13, -5, -35, -15, 4, 20, -24, -10, -11, -29, 48, 23, 4, -32, -7, 30, -11, -6),
    (15, -9, -12, -34, 22, -7, -44, -67, -28, 36, -55, -38, 6, -9, -21, -2, 24, 54, -56, 16, 3, -4, 0, 17, -30, 14, -6, 5, -19, 15, -23, -5, -43, 21, 10, -49, -11, -37, 9, -19, -10, 5, -11, -43, 6, -51, -23, -9, 5, 63, -51, 41, 10, -37, 34, 23, -23, 19, -43, 21, -39, 13, 22, 3, -11, -1, -9, -21, -15, 12, -35, -11, -21, 37, 10, -31, -12, -38, -3, -15, 19, 45, -28, -12, 35, -44, -17, 35, 2, 8, -33, -15, 2, -16, 26, -23, -35, 48, 29, -24, -3, -7, -10, 22, -1, 59, 6, -21, 3, -29, -34, -18, -9, -3, -52, -5, 18, -28, 29, 6, -16, -2, -25, -5, 17, -23, 5, -23, -27, 7, 30, -13, -21, -15, 7, -7, 19, 43, -44, -26, 1, 30, -32, -2, 32, -10, -10, 6, -6, -31, 24, 53, -32, -9, -24, 20, -13, 37, 43, 29, -19, -32, 22, -16, -13, -8, -1, -45, 22, 10, -52, -23, 31, 12, 10, 9, 6, 47, -5, -20, 13, -40, 42, 39, -11, -2, -23, 5, -17, 17, -36, -8, 1, -10, -18, -54, -34, 6, -30, -15, -41, 23, -3, 17, -36, 35, -15, -13, 0, 17, 7, 28, 21, -28, -2, -21, 1, -4, -48, -15, 5, -4, -13, 18, -20, -17, 24, -38, -19, -5, -8, 24, 42, 28, -5, 28, 17, 16, -5, -41, -15, 38, -14, 34, -16, -36, 25, 0, 7, 0, -32, -48, 28, -25, 0, 3, -16, -23, -38, -14, 40, 19, -36, 17, -7, 17, 16, -28, -9, 20, -38, -15, 1, -20, -18, 14, -30, -41, 36, -32, 14, -20, -39, -23, -6, 36, 0, -42, -11),
    (-28, -44, -30, -24, 22, 19, -19, 35, 14, -33, -43, 4, -26, -33, 12, -4, -9, -30, -45, -2, 5, -17, -6, 8, 16, 2, 2, 4, 16, -41, 5, -45, -20, 7, -38, 0, -11, 19, 37, 24, 43, -44, 9, -11, -47, 34, -35, -5, -33, -47, 36, -39, -17, -49, -38, -4, 17, -12, -41, 31, -24, 14, 6, -13, 21, -42, 9, 0, -2, -14, -1, -25, 11, 15, 37, -5, 31, 39, 18, -15, -12, 16, -35, -45, 18, -12, -52, -21, -25, 27, 32, 30, -34, 2, 13, 8, 37, -20, -21, -24, -1, 23, 6, 35, 19, 9, -29, 7, 9, -34, 2, 1, 17, 2, 12, 7, -9, -33, -8, 0, 28, 16, 33, -9, -11, -33, 53, 27, 23, -7, 29, 35, 24, 12, 29, -18, 8, -9, 7, -30, -10, 9, -8, 11, -24, 43, -18, -2, 28, 26, -15, 39, 29, 15, -10, 74, -5, 66, -13, 40, -6, -4, 15, 35, 4, -4, -23, -2, 7, -16, -20, 3, -18, 13, 57, 14, 5, 41, -88, 27, 32, 48, 22, 27, 34, -25, 2, 39, 4, 28, -42, 16, -5, 12, -21, -1, -16, 5, -19, 37, 27, 22, 15, -7, -21, -32, -23, -9, -60, 24, -36, 3, -18, -4, -6, 30, -30, 20, 9, 24, -24, -20, -14, 35, -15, -14, 31, 42, -37, -11, -45, -34, 9, -22, -8, 20, -31, -6, 11, -10, -24, -14, -19, 10, 19, -18, 46, -7, -41, 22, 27, -4, -27, 21, -5, 5, -17, -9, -35, 15, -48, -29, 8, -32, -19, -18, -27, 10, 1, -38, 30, 2, -21, -39, -3, -42, 8, -27, -4, -10, -34, 10, 0, -19, 19, 1, -35, -22, 0),
    (47, -17, 44, 14, 44, 2, 28, -1, 16, 6, 24, 21, -8, 16, -9, 18, -16, 6, -22, -12, 11, 14, -20, 44, -9, 35, 32, -36, 5, 1, 0, -29, 34, -14, 18, -52, 32, -3, -4, -15, -27, -23, -8, 5, 1, 15, 23, -12, -20, 12, 35, -15, -24, 21, 11, 28, -9, -35, 17, 15, -49, 47, -9, 26, -9, -6, 38, 33, 23, 10, 37, -16, -42, 2, -22, -46, 12, -10, 6, -7, -12, 7, 23, -45, -24, 19, 26, -15, 4, -15, 18, -46, -16, -2, 9, 7, -25, -10, -40, -26, -4, 13, 10, -66, 3, -25, -45, -21, 30, -10, 27, -6, 44, -33, -22, -39, 11, 23, 16, 8, 25, 4, -34, 16, -14, 43, 6, 8, -41, -24, -28, 2, 9, -5, -5, -30, -3, -15, -35, 1, -45, 8, 2, 2, -45, -50, 33, -10, -58, 9, 10, -27, -6, -44, -40, -26, -4, -6, 38, -9, -19, 29, -21, 45, -50, 25, 41, 24, -24, 20, -2, 7, 16, -9, -2, -40, -36, -28, 34, -37, 7, 5, 46, 5, -3, -1, -25, 7, 12, -3, 15, 8, -10, -25, -31, -26, -40, 7, -7, -26, -36, 3, -17, 18, 13, 23, 13, 12, -7, -13, 37, -30, -32, -38, -17, -2, 9, -19, -28, 16, -20, -32, 45, 36, 21, 24, 24, 7, -55, 24, 52, 8, 28, -5, -13, -8, -32, 28, -8, 24, -42, -6, 27, -17, 25, 15, -13, 27, 6, 18, -26, 6, -11, -14, -10, 23, -32, -15, -3, 7, 25, 31, -21, 26, 42, 7, 32, -13, -13, -43, 26, -14, -10, 13, -3, 31, 46, 26, 33, -8, -21, -7, 20, 43, 41, -7, -13, -27, -2),
    (-36, 28, -31, -34, -15, -42, -46, -39, 23, 18, -43, 45, 21, 27, -18, 1, 6, 20, -16, 34, 13, -27, -29, 2, 0, 15, -14, 5, 15, 10, -9, 14, -22, -27, -31, 24, 6, 33, 16, -13, 20, -6, -9, 6, 35, 23, -21, -24, -13, 27, 63, -35, -21, 40, 14, -15, 20, -15, -22, 18, -33, 23, 59, 8, -44, -35, -14, -20, -8, 7, -27, -38, -19, 32, -29, 20, -13, 20, -6, -15, 21, 25, 22, -28, -26, 25, -19, 15, 54, 3, -53, 7, -5, -27, 26, 14, -34, -3, -8, -48, 18, -31, 12, -52, -18, 20, -15, -12, 17, 8, -12, -13, -36, -52, 30, -6, 0, -21, -52, -9, -7, -30, 25, 14, -20, 9, 2, -41, -23, -11, -51, -6, -6, 27, -25, 7, 5, 16, -13, -36, -13, -26, -13, -32, -56, -27, 80, 7, -48, -19, -34, 11, -12, 3, -11, -19, -30, -6, 10, 35, 13, 9, -1, 10, -42, 2, 30, 15, 33, 28, 28, -25, -4, -9, 17, -16, -20, 15, 19, 3, 29, -13, -40, 1, 20, 47, 22, 17, -24, 1, -49, 11, -24, -23, -25, -14, 24, 5, 1, 3, -51, -36, 29, -18, 4, 10, -45, 28, 7, -13, 4, -11, -44, -7, 3, -8, 0, -22, -29, 27, 10, 31, 2, 0, -23, -2, 12, -19, -33, 14, 8, -31, 4, -1, -23, -35, 41, -43, -27, 42, 14, -30, 30, 46, -10, -4, -23, -32, -20, -7, 23, -20, -25, -28, 26, 34, 27, 16, 2, 34, -21, 39, -12, 11, 21, -12, 35, -46, 9, -40, 5, 29, 1, 10, -56, -34, 39, -36, -22, 25, 14, 11, 40, -18, -26, -1, -12, 24, -11),
    (16, 33, -20, -10, -29, 10, 21, 19, 14, 23, 14, -8, -39, 28, -6, -8, -32, -12, 24, 13, -45, -20, -10, -41, -9, -4, -16, -33, -7, 29, 38, 26, -30, -30, -2, 39, -19, -19, 29, -20, -18, -15, -7, -18, -30, 30, 30, -24, -27, 1, 19, -2, -5, 0, 23, 6, 26, 8, -5, -33, -45, -25, 37, 18, -48, -12, -17, -16, -3, 39, -1, 10, 25, 11, -2, -43, -28, -11, -54, -24, -8, -24, 12, -5, 31, 4, 11, 20, -12, 19, -13, -6, -13, 9, 8, -4, -25, -44, -17, -62, -7, -14, 46, -44, -14, -34, 3, 11, -51, -32, 6, 3, -40, -61, -32, -43, -15, -21, -38, -12, 8, -21, 46, 25, 0, 18, -16, 0, -5, 8, -14, 1, -12, -29, 38, 50, 8, 11, 15, -28, -28, 28, 36, -10, 18, -20, -14, -15, -20, 5, 11, -3, -30, -27, 35, 34, 18, 39, -17, 25, 5, 3, 2, -12, 31, 21, 43, -10, -10, 0, 41, -33, 13, 41, 37, -28, 44, 25, -50, -24, -22, 21, 15, 6, -35, 37, 27, 36, 13, 31, 28, 28, 20, -37, -10, 24, -15, 43, -10, 2, 9, 38, 4, 21, -20, 37, 8, 8, 8, 3, 6, 5, 26, -1, 3, -16, 11, -34, 14, -4, -21, -11, 36, -22, 31, -46, 15, 17, -17, 22, 39, -50, -36, -40, 36, 6, -24, 45, -11, -3, -18, -2, 22, 3, 6, -33, 29, -3, 57, -7, 17, -35, -37, 10, 10, -1, -1, 11, 20, -18, -28, -6, -24, -49, 11, -16, 26, 11, -38, -17, -13, -21, -44, 0, 14, 15, -15, -6, 30, 21, 35, -2, -16, 8, -5, -12, 20, -13, 6),
    (-14, -5, 18, 13, 2, -24, 30, 0, -45, -9, 6, -20, -30, -11, -88, -9, -26, -3, 1, 20, -27, -32, 26, -1, 6, 4, -30, 5, -47, -31, 3, 16, 17, 28, -21, -22, -6, -18, 23, -1, -24, 7, 8, -26, 8, -34, -77, 0, -54, 17, -12, 27, -24, 11, -1, 19, -16, -36, -2, 35, -41, -44, -14, 14, 18, 22, 2, -8, 21, 25, -33, 5, -42, -19, -11, -33, 1, -36, -65, 9, -44, 22, -32, 18, 13, 17, 33, -18, -9, -27, -8, -19, -44, -3, 32, -2, 27, 8, 47, 27, 14, -23, -14, 34, 31, 13, -4, 17, 5, -17, 65, -5, 24, -37, 15, 23, 10, 0, 31, -19, -19, 5, 31, -5, 12, 52, -21, -15, -13, -11, 24, 35, 32, -25, -11, -5, 22, 35, -33, 6, 38, 8, 60, 19, 35, 20, -6, 27, -13, -22, 35, 7, -9, 36, 20, 11, 7, 28, 0, -21, 29, 6, 24, 6, -9, -8, 37, 15, 5, 17, 21, 6, 27, 13, 31, -16, 9, -19, -32, 8, 11, -51, 16, -26, -6, 31, 10, 10, 1, 1, 21, 3, -11, -21, -3, 25, -7, -1, -13, -3, -1, -40, -34, 28, -17, -7, 22, 13, 36, 11, 2, -11, -31, -24, -71, -27, -2, -6, -3, -32, 18, 4, -4, -7, 6, 26, -39, 28, 15, 12, -15, -29, -33, -27, -7, 22, -32, 13, 14, -34, -16, -31, 23, 2, -8, -8, -56, -37, -14, -14, 1, -37, -16, -5, 19, -40, -11, 24, -36, 42, 39, -29, -39, 32, 1, 20, -8, 17, -1, -4, -13, -47, -18, -21, -21, -29, -2, 5, -59, -20, -12, 3, -16, 6, 24, 8, -16, -51, -7),
    (4, -11, -2, -46, -44, -16, 19, 27, -51, -43, -42, -51, -4, -36, -39, 9, 3, 0, -57, -2, -38, -2, 26, 9, 3, 7, -15, -11, -68, 19, 25, -57, -2, -29, -32, -22, -47, -22, 7, -16, 16, -9, -52, 5, 28, -15, -14, 9, 3, 19, -1, 16, -24, 31, -54, 1, -57, 6, -17, -22, 11, -28, 6, 17, -14, 0, 10, -23, 12, -39, -55, -9, 5, -26, 15, 7, -18, -12, -6, 59, 27, -20, 3, -4, -21, 27, -63, 15, 10, 27, 23, 5, 29, -14, -15, 38, -9, 28, 9, -31, -8, 13, 17, -27, 5, 27, -7, -14, -9, 35, 48, -6, 25, 45, -13, 39, 34, -7, 11, -4, 19, -2, 3, -9, -22, 24, 8, 24, -11, 12, 17, -38, 4, -26, 35, -36, 11, 6, 26, -38, -1, -14, 31, 27, 1, 32, -59, 17, 1, 44, 19, -16, 0, 12, 21, -14, -13, -5, 54, -13, 9, -6, 27, -45, -24, 2, 13, -39, -10, 31, -32, 10, 5, -17, 12, 38, 9, 22, -5, 22, -17, 12, -52, 9, -4, -5, -2, 6, -22, -8, -31, 26, -35, -12, -93, -23, -42, 10, -26, 12, 1, -28, -16, 6, -35, -22, 5, -17, -32, -2, 40, -6, -63, -9, -42, -61, 13, 17, -13, -34, 11, -30, 28, 15, 15, -23, -25, 36, 14, -11, 12, 25, -9, 36, 4, -12, 27, -39, 26, -9, 25, 9, -45, -21, 3, -15, -3, 13, 22, 9, 26, -34, 10, -35, 12, -19, -9, -21, 18, 6, 16, -24, -18, 29, 12, 2, -9, -8, 8, -45, 4, 19, 10, 1, -42, -15, -42, -19, -66, 23, -38, 26, 16, -41, -13, 49, -31, -34, -7),
    (32, -51, -18, -26, 18, 47, -14, 26, -18, -5, -20, 1, -47, 44, 32, 31, -38, -32, 9, -17, -28, -27, -29, -27, -5, -24, -49, -1, -8, 26, 34, 37, -48, 12, 14, 8, -53, 11, -3, 13, 4, 28, -12, 32, -11, 8, 48, -28, 32, -23, 5, -15, -7, -37, -21, -8, -19, -11, -7, -20, -13, 22, 42, -3, -47, 4, 1, -22, -9, -60, 35, 1, 21, -18, -45, 9, -39, -17, -5, -4, 34, -56, -3, 25, 33, 40, -7, -21, 36, 22, 8, -2, 67, -4, -15, -23, 26, 4, -40, -15, -9, 21, 49, 15, -9, -1, -3, 0, -6, 31, 27, 33, -12, 10, -3, -15, -16, 6, 31, 22, -16, -35, -38, 36, -23, 45, -48, 22, -15, 24, -36, -5, -7, 15, 14, 21, 0, -8, -9, -6, -32, 41, 1, -48, 36, -36, 22, -4, -3, 17, 4, 39, -22, 23, -17, -13, -4, 41, -31, -48, 7, -33, -12, 47, 54, -3, 26, 33, -50, 26, -20, -34, 21, 1, -16, -59, 38, 8, 17, -7, -7, 19, 13, 26, 21, 26, 17, 21, 24, 17, 1, -38, -29, -2, -19, -9, -53, 9, 8, -4, 26, -32, 21, -17, 7, -7, 10, -23, -41, -19, -3, -20, 26, -12, 16, 17, -10, 9, 23, 24, 9, 8, -7, -5, 3, 0, 20, -3, -31, -34, -7, -2, 33, -36, 8, -32, -37, 18, -18, 19, -22, 21, -30, 28, -22, 1, 33, 3, -8, -21, -39, -13, 17, -9, 49, -16, 2, -39, 9, 16, 2, 17, 18, 5, 6, -34, 27, -20, 24, -19, 32, -24, 10, 46, 15, -40, -18, 2, -15, 4, 7, -18, -43, -40, -14, -5, 27, -16, 7)
  );
  ----------------
  CONSTANT Layer_7_Columns    : NATURAL := 8;
  CONSTANT Layer_7_Rows       : NATURAL := 8;
  CONSTANT Layer_7_Strides    : NATURAL := 2;
  CONSTANT Layer_7_Activation : Activation_T := relu;
  CONSTANT Layer_7_Padding    : Padding_T := same;
  CONSTANT Layer_7_Values     : NATURAL := 32;
  CONSTANT Layer_7_Filter_X   : NATURAL := 3;
  CONSTANT Layer_7_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_7_Filters    : NATURAL := 48;
  CONSTANT Layer_7_Inputs     : NATURAL := 289;
  CONSTANT Layer_7_Out_Offset : INTEGER := 3;
  CONSTANT Layer_7_Offset     : INTEGER := -1;
  CONSTANT Layer_7 : CNN_Weights_T(0 to Layer_7_Filters-1, 0 to Layer_7_Inputs-1) :=
  (
    (-22, -17, -1, 4, -3, -9, -22, 2, -11, -20, -12, -3, -42, 37, 27, 16, 28, 22, -1, -17, 2, -4, -49, -6, 15, -17, -42, -28, -54, -18, 14, -31, -46, -1, -13, -18, -21, -21, -8, 30, 17, -22, 13, 13, -27, -13, 6, 19, 3, 18, 45, -27, -3, 36, -22, 21, 24, -16, -33, -31, -29, -10, -20, -21, -22, -14, 28, -18, 6, 14, 10, -36, -1, -7, 33, -31, -33, 1, 6, -31, -6, 16, -28, -36, 50, 40, 25, -1, 15, 24, 26, -16, -9, -17, 18, 18, 7, 28, 13, -11, 16, 10, -3, -15, 37, 40, 41, -25, -12, -15, -3, 40, 30, 5, 3, 4, -30, 5, -49, -18, 45, -25, -26, -5, -35, -33, -1, -30, -3, 39, -2, -12, 5, 25, 22, -10, -21, 33, -35, -19, 4, 35, -22, -2, -1, -31, 29, -25, -23, -19, -35, -8, 34, -50, -14, 2, -35, -39, 34, -12, 20, 41, -25, -7, -31, 36, 11, -26, 9, 25, -18, 14, -18, 49, -4, 7, 12, -42, 14, -24, -12, 36, 13, 24, 11, -42, -16, -21, -20, -28, 53, -12, 29, -47, -15, -10, -15, -8, -26, 0, 3, 27, -26, 16, -3, 28, 6, 12, 23, -35, 17, -21, 27, 12, -10, -9, 43, -26, -2, -16, -10, -21, 30, -32, 39, -19, 36, 7, -6, 36, 4, 32, -3, 30, -12, -8, 25, 26, -26, 54, 32, -49, 8, 16, 9, 24, -12, -6, 37, -28, -9, 3, -11, -13, 31, -34, 37, 17, 28, 6, 9, 27, -22, 4, -19, 29, -29, 0, 36, 23, -9, 18, -28, -26, 2, -22, 18, 20, -6, -6, 41, -5, -36, -26, -14, -1, 33, 50, -9),
    (-9, -16, -15, 40, 38, -53, -26, -7, -16, 1, -12, 3, 25, -50, -5, -7, 22, 41, -34, 13, 26, 14, 8, 10, 24, 29, -9, -10, -4, 45, -34, 20, 35, 0, -11, 18, 25, -47, -8, 21, 20, -36, -33, 42, 45, -54, 16, -23, 24, 10, 0, 23, -27, -27, -10, 29, -11, 25, -5, 5, 25, 0, -26, -17, 34, -25, 11, 30, -23, 1, -6, 44, 10, -58, 5, 9, -15, -16, 12, -29, 40, -23, -28, 34, -6, -11, 8, 31, 14, 17, 21, -3, -15, 10, -28, 12, 8, 3, 7, -40, -9, -24, -20, 34, 18, -4, -1, -27, -14, -65, 51, 6, -14, 10, -27, 22, -14, 6, -5, 25, -15, 20, 6, 15, -45, 14, -19, -20, -13, -23, 31, 1, -19, -45, 18, 53, 19, -33, 21, 9, -17, 16, 48, -42, -2, 51, -60, 32, -37, -10, -7, -4, -24, 29, 20, 17, -16, 7, -74, -50, 38, -6, -12, -1, -38, -6, -20, 0, 46, -31, -16, 0, 39, 0, 4, -2, -5, 27, -26, -3, 14, -36, 17, -17, 8, 39, 32, 10, 31, 8, -65, 15, -43, 18, -3, -29, -12, 5, -21, -9, -29, -23, -4, 0, 6, 3, 23, -11, 16, 3, 2, -7, -36, -47, 22, 19, -9, -6, -23, -6, 9, -12, -25, 5, 34, -23, 8, -56, -53, -29, -23, -8, -34, -27, -11, -42, -17, -35, 42, 5, -2, 30, -6, -29, -38, -42, 36, -1, -44, -45, 16, 39, 3, 26, -70, -11, -13, -40, -55, -9, -31, -8, -43, 4, -31, -24, 25, 3, 23, 3, 15, 46, 13, 23, -16, 60, -42, -23, 18, 25, -8, 37, 40, 28, 21, 18, -56, 0, 47),
    (39, 14, -42, 8, 25, -12, -26, -12, -20, -17, 31, -51, -27, -20, -13, -33, 3, 8, 37, -18, 18, -35, 17, 3, -15, -3, -17, -17, -36, 1, -39, -12, 28, 26, -27, -7, 29, -28, -21, 1, 32, 20, 56, -26, 23, -19, -29, -33, -19, 12, 12, -10, -29, -23, 33, 7, -6, -19, -61, -30, 4, 31, -40, -39, -7, -9, -8, -1, 34, -14, 21, 4, 24, -28, 8, 17, 25, 2, -55, 1, -12, 10, -13, -2, -34, -11, 7, -11, -25, -3, -35, -14, 24, 47, 6, -22, 26, 4, -56, 20, -2, 17, -11, 7, -9, -18, 22, -20, -38, -12, -21, -41, 11, 50, -16, 10, -25, -49, 29, 41, 15, 13, 12, -28, 27, 47, 22, -9, 21, 35, -66, 45, 53, -44, -34, -3, -16, -20, 52, -2, 24, 8, 5, -46, 39, 46, 5, -25, -1, -53, -1, 18, -17, 0, 1, 1, -15, 44, 15, -19, 10, 17, -25, 18, 31, -1, -18, 4, -27, -33, 30, -2, 17, -5, -1, -30, 28, -32, 11, -43, -41, -4, 31, 14, -26, -46, -6, -5, -7, 18, -9, -23, 32, 0, -7, 25, 26, -2, -21, 27, 27, -27, 3, -15, -1, 12, -17, 12, 11, 45, -24, -6, 34, -10, 25, -3, -5, 2, 9, -15, 10, 36, 14, 34, -29, 33, -12, 43, 37, 51, -24, -3, -4, -44, -7, -21, 38, -8, 8, -16, -9, 29, -6, 12, 23, -19, 1, 7, -44, 2, -2, 2, -11, 32, 28, -3, 33, 12, -15, 1, 13, 36, -28, 20, -24, -25, -9, 17, 1, -40, -29, -47, -4, -18, -8, 1, -32, 7, 26, -23, -2, -29, 3, -21, -12, 14, 26, -8, 11),
    (-28, -22, 26, -21, -20, -3, -4, 13, 0, -25, 1, -23, -4, -8, 58, -21, 59, 26, 2, -18, 1, -41, 1, 2, 24, 12, -63, -27, -6, -23, -2, -7, -34, -49, -38, 3, 34, 2, -29, 12, 5, -45, 61, -11, 28, 26, 61, -6, 51, 30, -31, -16, -38, -25, -14, 8, -27, -12, 6, -43, -17, -23, 15, 31, 6, -42, -18, 24, 23, -20, -36, 1, 14, -6, 32, -12, -32, -4, 37, 19, -4, 52, -9, -9, -2, -9, -18, 8, -10, 9, -23, 16, 19, 0, -26, 8, -33, -36, 20, -13, 10, 7, -19, 20, 55, -52, 12, -12, -12, 18, 68, 6, 46, 13, 7, 7, -40, -16, 0, -22, -50, -19, -18, -37, 7, -27, 3, -4, -31, -31, -18, -11, 1, 18, 8, 23, 27, -63, 42, -21, -27, 2, 58, -11, 22, 52, -26, -8, 5, -5, 3, 18, -19, -2, 2, -40, -35, -1, 24, 14, 5, -39, -58, 11, 49, -14, -6, 36, 10, -22, 54, -13, 11, -13, 31, 23, -9, 24, 10, 20, 16, -16, -20, -1, -16, 17, -11, -42, 12, 34, 11, -22, -37, -15, -39, 5, 14, 6, 31, 1, 9, -18, 54, -3, 3, -25, 28, -19, 5, 32, 5, 30, 12, -53, 6, -7, -29, -35, 9, 17, -15, 3, -7, -3, -4, -34, 12, -7, 2, 13, -26, 8, 16, -5, 7, -8, -9, 20, 44, -8, -13, 3, 32, 9, 26, -19, -17, -2, 9, -26, -16, 19, -18, 21, -10, 16, 16, 5, -17, 14, 26, 20, 31, -6, 1, 18, -7, 10, -29, 3, -39, -32, -14, -1, -1, -20, 25, 21, -8, 38, 31, -9, 37, -36, 10, 9, -11, -13, 11),
    (-22, 40, -13, -37, -9, -4, -38, -61, -9, -13, -36, -13, 24, 24, -3, -9, 30, 19, -40, 5, 18, 10, 18, -14, -13, 19, -2, 24, 23, -24, 7, 12, -34, -2, 31, 0, 0, -1, 2, -55, 10, 6, -33, -17, 22, -19, -23, -14, 20, -9, -15, 49, -16, 8, -19, -6, -6, 28, -40, 6, 11, -41, 4, -26, 2, 3, -7, -15, -30, 25, 31, 5, 26, -43, 6, -7, -13, -41, -30, -12, -2, 20, -23, -10, 32, -21, -2, -2, -5, 34, 13, -6, 9, -9, 4, -13, -32, 41, 21, -26, 9, -9, 8, -22, 19, 32, 9, -29, -17, -23, -20, 26, -23, 10, 1, 15, -38, 35, 6, 12, -6, 24, 5, -34, -4, -9, -2, 1, -29, 59, 24, -7, -5, -9, 17, 23, 2, -7, -8, 1, -20, -36, 23, 4, -17, 44, -33, 16, 40, 27, -6, 21, 3, 17, -37, 34, 26, 6, -25, 1, 15, 1, -26, 13, -4, -39, -22, -38, -21, -12, -25, -1, -1, -19, 9, 19, -1, 38, -46, -1, 31, 2, -3, 28, 22, 20, -2, 26, 22, 37, -40, -47, -43, 55, -26, 31, 23, -37, 41, 6, -4, 16, 0, 4, 7, -18, -16, 30, -16, -16, 10, -29, -24, 36, -5, 9, -10, 4, 28, -8, 29, 17, 15, 8, -11, 26, 33, 3, -33, -16, 5, -32, -27, 28, 6, -31, -39, -21, -21, 1, 4, 20, -12, -29, -21, -14, 12, -35, -20, 30, -13, 4, 7, 23, 18, -1, 19, 5, 23, 32, 20, 26, 17, -4, -34, 10, 13, 0, 19, 10, -31, -2, -26, 11, -16, -8, -20, 11, -2, 2, 29, 7, 36, -8, 31, -17, -35, 35, -11),
    (-35, 6, 13, 12, 25, -14, -26, 34, -33, -33, -4, -12, -10, -19, -3, -37, 13, 7, -36, 12, 1, -38, -16, 25, -48, 6, -16, 24, 15, 13, 19, 68, -44, -13, 3, 12, 17, -33, -20, 49, -7, -40, -3, -24, -25, 20, -47, -28, 9, -16, -7, 1, -19, -18, -20, -17, -14, -2, 12, -21, 46, -21, 0, 46, -41, -8, 7, -16, 10, -11, -33, 1, 1, 18, -16, 26, 14, 16, -11, -20, 37, -44, 12, 8, -19, -33, 9, 11, -10, 12, -29, -7, 34, 3, -47, 7, -5, 7, -39, 19, 44, 19, -54, 27, -36, -4, 18, 31, 4, -14, -24, 17, 7, 28, -48, 15, 8, 18, 25, -23, -10, -42, -27, -18, 1, 40, 12, 1, 24, -31, 0, 0, 29, -39, -70, 40, -36, -26, 40, -26, -43, -11, -3, 8, 17, 2, 15, 31, -4, -2, -19, -26, 2, -46, -5, -36, -39, 51, -5, -4, 2, -16, 6, 21, 23, 3, -35, 45, -9, -8, 7, 26, 26, -5, -42, -34, 9, 5, -16, 1, -37, 7, -34, 0, -10, -1, 45, -20, -4, 13, -41, -12, 32, 19, 30, 8, 28, 1, 19, -16, -6, 27, 13, 21, -4, -12, -3, 10, -38, 25, 2, -16, -17, 37, 6, 34, 16, -6, -11, 22, -29, 26, -2, -52, 32, 26, -3, 29, 40, 1, -1, -14, -7, -24, -1, 6, -14, -19, -46, 1, -28, 33, -4, -36, 3, -30, 3, 24, -24, -2, -28, 12, -25, -20, -6, -39, -11, 47, -10, 28, 1, -10, -13, 25, 34, -35, 18, -15, 28, -40, -1, 11, 0, -11, 34, 9, -19, -55, -14, 40, -11, -11, -2, 20, -26, -40, 0, 23, -8),
    (17, -3, -15, -11, 25, 30, -24, -14, 19, -11, 22, -40, 0, -35, -20, 9, -3, 27, -36, 22, 21, 7, -24, 26, 17, 5, 19, 40, -16, 22, 29, -43, -24, 11, -30, 8, 27, 53, -24, 20, 15, 20, 6, -14, -9, 25, -40, 41, -3, 50, 19, -12, 34, -1, -22, 22, 36, -5, -7, 25, -35, 28, 29, -55, -2, 19, 24, -43, -22, 8, 0, 11, 8, 13, -13, -4, -9, 32, 0, -8, -14, 32, -4, 28, -2, -10, 9, 3, -3, -18, -6, -13, 13, 19, 55, -31, -8, 4, 19, 21, 30, -15, 1, -18, 14, 17, -15, -5, -26, 36, -36, 13, -23, -15, -10, 23, -9, -20, -21, 14, 11, -23, 2, 23, 3, 38, 23, 2, 12, 15, -14, -11, -22, 33, -2, 19, -4, -9, 5, -53, 39, 21, -53, 42, 20, 65, -5, -7, 32, -31, -11, 19, 26, -4, 18, 33, 19, 39, 57, -42, -24, 3, -26, -18, -43, 36, 5, 8, 2, 10, 2, 16, -11, 60, -37, 32, -11, 44, 9, -27, -13, -28, -11, -7, 34, -23, 9, -22, 31, 2, 54, -13, -20, -8, 6, 27, 20, 20, 9, -39, 25, -15, 19, -29, -46, -2, -8, 17, -5, -27, 1, -9, -8, -31, -4, 31, -20, -2, 9, 16, -6, 11, -7, 16, 10, -40, 5, 21, -19, 3, -2, -4, -24, -1, -9, -2, -1, 6, -27, 7, -30, 20, -7, 35, 18, 29, -5, -7, -26, 6, 34, 37, -22, 28, 12, 21, -26, -11, 3, 40, 11, 4, -30, -26, -43, -6, -16, -55, -16, 37, 5, -12, 27, 2, -24, 16, -31, -13, -24, -18, 27, 6, -23, 45, 23, -16, -10, 29, -13),
    (-7, 6, 2, -46, -17, 21, -8, -4, 17, -11, 19, 2, 28, -20, 36, 27, 7, 41, -31, 8, 12, -49, 2, 44, 19, 7, -19, -2, 6, -47, 15, -34, 35, 29, -34, -21, -22, 4, 29, -2, 48, -20, -18, 11, 15, 1, 33, 47, -23, 42, -42, 50, 5, -38, -10, 30, -9, 31, 21, -14, 13, -8, -27, 2, 16, -1, -36, -23, -12, 2, 28, -20, 18, -6, 17, 3, -22, -6, 4, 27, -33, 4, -31, 30, -13, 24, 7, 10, -17, 23, -16, -30, 4, -3, 10, -38, 33, -1, 8, -8, -11, -30, -29, -6, 14, -9, 9, -22, -18, 5, 45, 31, 19, 5, -41, 28, -9, -70, -2, 43, -39, 14, -15, 14, -25, -31, -32, -22, -10, 19, 4, -8, -32, -31, 26, -21, -12, 7, -14, 1, 42, -12, 20, 15, -17, 50, -29, 4, -13, -71, -19, 43, 3, 6, 32, -7, -27, -34, -11, -26, -26, -15, -1, 13, 25, 5, 6, 26, 3, 25, 27, -27, 22, 10, 43, 13, -11, 57, -64, 39, 0, -13, 12, -12, 25, 22, 19, -11, -8, 30, 19, -28, 13, -22, -22, 1, 4, 32, -13, 5, 12, 8, -12, -1, -27, -40, 40, -3, 25, 10, -13, 40, -41, -54, -15, 19, -47, 32, -15, 9, -38, -3, -32, 5, -6, -8, -15, -34, 19, 17, -19, 1, 0, -35, -10, 9, 15, -41, 5, -28, 27, 27, -21, 32, -41, -53, 4, 20, -33, -1, 28, -7, -7, -27, -22, -11, 4, -18, -27, -49, -25, 16, -37, -33, 27, -18, -17, -4, -3, -8, 27, -44, -18, 29, 8, 18, -54, -48, 40, 24, -15, 39, 21, 44, -35, -5, -26, 25, 9),
    (11, -10, -27, 27, 25, 25, -2, 53, -6, 24, 15, -30, 6, -51, 38, 26, -21, 14, 13, 13, -41, 22, -39, -3, -38, 25, -36, 10, 16, -5, 27, -48, 37, -3, -18, 12, 10, 57, -8, -8, -28, 26, 27, 15, -35, -33, 33, 58, -36, -4, 2, -8, -13, 3, 7, 7, 17, 21, 6, 34, -41, -47, -1, -47, 38, 33, -4, -7, 5, 18, -17, 21, 6, -39, 13, 0, -12, -22, 7, 1, -20, 18, -39, -23, -21, 6, -4, -1, 32, 36, -17, -21, -12, -47, -8, -24, 19, -44, -49, 9, 11, 3, -23, 3, 17, -36, -24, -27, 26, -43, -12, 47, -1, -10, -25, 0, -2, 10, -15, 42, 38, 56, 23, 38, 2, -31, 3, 21, 29, -41, -24, -12, 2, 16, 6, 40, 41, -12, -6, -31, -3, 14, -3, 18, -16, -17, -1, 26, 22, -4, -32, 7, -10, 39, -18, 1, 29, 43, 5, 22, 22, 3, -8, 6, 18, 51, 23, 27, -21, 34, -21, -3, 23, -24, 13, 33, -21, 5, 20, -14, 26, -42, -11, 50, 25, -12, 33, 24, -13, -10, -10, -13, -1, -59, -18, 2, 37, -10, -31, -38, -42, 15, -15, 1, -6, 27, -43, 18, -35, 1, -1, 32, 32, -1, -16, -19, 6, 14, 20, -4, 19, 48, 0, 50, -8, -46, 2, -8, 32, -11, 26, -37, 5, 16, -24, -13, 15, 0, -33, 23, -21, -20, 15, 2, -2, -20, -6, 7, -1, -1, 44, 23, -26, 22, -26, 20, 21, 20, -27, -25, 36, 19, 5, -31, 7, -23, -36, 0, 37, -22, 13, 19, 1, 12, -29, -11, 27, -6, 6, 13, -13, 3, 29, 36, -24, 28, -19, -14, -10),
    (-22, -23, -13, 30, 1, -34, -12, 39, -1, 1, 15, 39, 7, -39, 1, -24, -8, 25, 2, 37, -22, -37, -9, 15, -52, -35, 19, -38, 15, 7, -33, 5, -4, -36, -60, 48, 38, 16, -38, -3, 13, 15, 30, 6, 1, -20, -26, -30, -17, 48, -20, -11, 26, -23, 35, 52, 12, -3, 10, -30, -23, 31, -38, 17, -20, -3, -55, 1, 49, 22, -30, 48, -38, -6, 36, -16, -2, -21, -2, 13, 18, 11, -5, -34, 25, -6, 2, 9, 28, -19, -23, -14, 13, 30, -12, -10, -12, -23, -55, 9, 41, 7, -21, 20, 11, -20, 1, -19, 34, -25, -22, -4, 30, 26, -24, 7, 21, -15, -10, 28, 2, -17, 10, -1, -50, 14, -1, 39, 13, 7, -16, 21, 31, 23, 7, 25, -4, 12, -1, -29, 3, 1, -28, 7, -6, 23, 15, 21, 3, -31, -21, 18, 27, 8, 42, -12, -57, 41, 2, 10, 21, -32, -7, 27, 1, 21, 34, -24, 27, -17, 37, 5, -6, -34, -17, 1, 14, 45, -27, -5, 11, -37, 25, 3, 2, -6, 37, 30, 20, 30, -25, -4, 11, -15, 6, -26, 20, 29, -5, 41, 29, -10, 13, 0, -17, -3, 12, 12, 19, 14, 7, -24, 17, -48, -32, 33, -7, 24, 10, -32, 9, 3, -8, -13, -15, 18, -17, -17, -44, 16, 40, 29, 15, -6, -15, -46, -16, -21, 9, 25, 27, 25, -5, -26, -17, -35, 6, 38, 4, 8, 30, -27, -14, -2, -12, -24, -21, 9, -6, -33, -73, 6, 28, -57, -28, -34, 10, -25, -24, 23, 26, -27, 20, 24, -21, -32, 3, -8, -7, -14, -48, -26, 20, -24, -8, -13, 31, -40, -1),
    (-12, -4, 28, 5, -20, 28, 2, -34, 42, 32, -2, -14, -26, -26, 0, -15, -48, -55, -1, -45, -20, 36, 30, 21, 48, 20, 20, 15, 29, -26, 34, -2, 13, 11, 39, 6, -36, 12, -27, -46, -16, 34, -1, 16, -13, 31, -5, -27, -21, -54, 11, -3, 28, 29, 38, 12, -5, 26, -18, 10, 27, 0, 12, 15, 8, -11, -3, -23, -3, 12, -45, -43, -29, 10, 23, 4, 7, -16, -39, -31, -36, 5, -13, 7, -5, -18, 20, 16, 40, -12, -26, 13, 18, 27, 9, -40, -6, 6, -13, -3, -12, 38, 13, 5, -6, 25, 2, -1, -18, 8, 11, -18, 31, -37, 10, -50, -23, 10, 12, 28, -26, 14, 20, -23, -9, -38, -25, -26, -25, -28, 40, -29, -19, 34, -5, -9, 22, 0, 0, 10, 14, 43, 60, -35, 24, -15, -22, 4, 15, 35, -28, -1, 17, -11, -35, 33, 62, -20, -6, -18, -42, -45, 31, -21, -45, 17, 11, -35, -22, -33, 28, 1, 20, 24, 36, -21, -1, -33, -26, -48, 4, 16, -17, 6, -24, 4, -34, 46, 20, -37, 14, 6, -4, -33, 24, -11, -24, 4, 9, 19, 12, -16, 7, -11, 34, 9, -5, -23, 29, -39, 6, 17, 10, 10, -1, 8, -11, -4, 54, -22, 54, 9, 6, 52, -1, -11, -10, 10, -27, -46, -3, 36, -20, -7, 15, -46, 38, -18, -19, 6, 16, -14, 10, 8, 19, -3, -26, -12, -38, 2, 35, -15, 43, 3, -36, 7, 12, 10, -26, -11, 7, 9, -12, 29, 9, 11, 21, -14, 56, -30, -12, 20, 29, -19, 10, 30, -39, -6, -31, -14, 0, -1, 2, 31, -1, 3, -49, 8, -6),
    (1, 22, 1, 16, -1, -6, -54, -18, -29, 45, 20, -29, -28, -14, 1, 42, -16, -30, 27, -27, -6, -23, -20, 6, -20, 17, 24, -15, 17, -19, -3, -1, 20, 38, -9, -4, 18, -20, 22, -3, 21, 24, -24, 2, 20, 13, 23, 16, -9, -6, -37, -14, -31, -15, -7, 42, 22, -1, 26, 35, -23, -29, -10, -34, 19, -43, 20, 19, 16, -12, -18, -31, 9, 27, 5, -6, -10, -27, -39, 10, -42, 4, -13, 7, 5, -25, -22, 2, 35, -27, 21, 11, 34, 2, 15, 5, 12, -1, 38, -28, -64, 3, -35, -10, 18, 34, -17, -3, 0, -30, -2, 37, 31, -45, -2, -21, -15, -3, -15, 24, -35, 20, 1, 37, -33, -54, 6, -64, -32, 45, 53, -21, -45, -6, -15, -32, 30, 24, -18, -43, 22, -26, -5, 4, 30, 8, -8, -12, -25, -30, -34, 37, -14, -12, -26, 50, -20, -25, 29, -40, -8, 22, 27, 22, -25, -1, -19, -41, 29, -6, -18, -20, -15, -10, 1, 15, -27, 4, 3, 3, 9, -22, -20, 20, 8, -14, 25, -3, -31, -21, 37, -47, 17, 17, 27, 35, -40, 1, -11, 13, 9, -18, -17, -24, 17, 5, 32, 8, 10, -2, 4, 16, 10, -49, -33, 28, 1, -34, -14, -17, -9, 14, 28, -37, -12, 7, 8, 7, -39, -31, -31, 4, 0, -25, -52, -34, -18, -30, 1, 36, -17, 27, -17, 15, -54, -18, -26, 39, 19, -20, -40, 30, -1, -9, 43, -27, 14, 3, 3, 25, -36, -26, 14, -29, 17, 12, 40, -45, -9, -30, -9, -16, -19, 31, 22, 23, 1, -42, -4, 21, 3, 27, 1, -5, -1, 19, 12, -32, -4),
    (-39, -25, -25, 9, 30, -6, -33, -39, 10, 37, -21, -33, -37, -41, -23, 19, 11, -18, -22, -36, -3, -28, 20, 19, 43, -19, -11, 18, -31, 32, 0, -4, -4, -25, -66, 11, 54, 11, -7, -17, 9, 53, 6, -27, -9, 16, -28, 10, 20, 1, -9, -34, -49, -18, 11, -12, -3, -18, -30, -13, 13, 10, 7, 19, 24, -10, -57, 24, -9, -24, 4, -2, 10, 25, -26, -7, 9, 18, -37, 1, 8, 31, -11, 0, -52, -12, -36, -11, 27, 22, -34, 40, 26, 27, -6, -5, 11, -4, -20, 29, 46, -37, 29, -25, 13, 22, 7, 30, -29, 46, -14, -40, 8, 16, 35, -2, -21, 34, 23, 13, 0, -21, -8, -30, -12, 56, -22, -12, 3, 5, 22, 22, 11, -41, 52, 23, 11, -1, -32, 28, -37, 27, -38, -17, 16, -11, 39, -22, 23, 14, 23, -26, -21, -31, 19, -33, -6, 16, 2, -27, 15, 16, -25, 22, -16, -68, 25, -13, 10, 14, -11, 48, 36, 2, 4, 22, 27, -24, 68, -20, -26, 10, -17, -1, -19, -11, 39, 40, -14, -34, -13, -31, 29, -10, 34, 15, 35, -45, 21, -22, -18, -4, 14, 43, 18, -31, 1, 2, -17, -14, -8, -19, -31, 51, 25, -21, -28, -3, 16, -66, 2, -16, -14, 18, -16, -20, 14, 36, -2, -22, -23, 13, -15, -15, -2, 47, -16, -24, -21, 6, -4, -74, 7, -15, 23, 11, 17, 9, -40, 9, 16, -8, 11, -4, -19, -21, -27, -31, 7, 31, 13, -28, -42, -26, -10, 4, -5, 32, 16, 4, -3, 4, 32, -8, -17, 1, -14, 9, -13, 20, -26, 8, -17, -25, 0, 9, 8, -23, 6),
    (12, 27, -45, 31, 12, -31, 27, 24, 6, 48, -8, 12, 7, -4, -27, 37, -26, 21, 39, -1, -25, 12, 30, -21, -39, 37, 0, 33, 38, -33, 12, -3, 45, 44, -49, 0, 2, -23, 31, 15, -13, -2, -2, 16, 33, 14, -19, 10, -12, 24, 39, 31, 18, 27, 50, 4, 7, 26, 40, 25, 4, -19, 17, 8, -21, 13, -2, -10, 19, -11, 6, -14, 2, -36, -18, 10, -26, 11, -1, -3, 2, 36, 34, -8, -10, 55, 14, 29, 4, 10, 33, 14, -23, -8, -18, -10, 32, -8, 48, -11, 2, 19, 28, 35, 36, 15, -45, 36, -5, 0, 1, 37, 1, -28, 15, 1, -19, 18, 17, 20, -35, 0, -6, 11, 46, 0, -25, -18, 12, -1, -10, 15, 30, -27, 14, -2, 8, -34, -31, 49, 20, -24, -51, 35, -28, -48, 49, -8, -20, 25, 26, 3, -22, 18, 30, 42, 35, -44, -12, -56, 32, 24, 0, 3, 15, 28, -3, 18, 9, -25, -25, 44, -15, -8, -36, 9, -13, -38, 24, -2, -22, 40, 24, 3, 14, 45, 21, 1, -13, -28, -22, 1, 4, -38, -31, -32, 13, -14, -12, -17, 32, 29, -53, -11, 13, -24, -1, 22, -5, -4, 25, 19, 4, 5, 3, 0, -6, 20, -2, -30, 21, -4, -2, -15, 16, -40, 8, 2, -13, 20, -36, -2, -15, 0, -4, 14, -36, -49, -5, 29, -14, -23, 43, 27, 22, -19, -15, -7, -4, 26, -47, -16, 39, -29, -15, -26, 11, -15, -7, -38, 33, 38, -3, 15, -23, -29, -36, 23, -14, -62, 16, 16, 15, -63, 12, 0, -13, -6, -47, -5, 2, -14, -27, 14, -20, -28, -12, -14, 9),
    (10, 14, -34, 3, -23, 7, 12, -1, 36, -10, 5, -10, 27, 9, -17, -10, 3, 13, 21, 48, 0, 12, -48, 5, 7, -1, 26, 35, -60, -14, 7, 23, 15, -4, -39, 34, 11, -1, 36, 6, 24, -50, 14, 16, -8, 20, 18, 2, 21, 2, -22, 25, -27, -19, -9, 21, -11, 27, 24, -21, -50, -1, 10, 24, -7, 21, -46, -53, -42, 46, -16, -35, 5, -5, 0, -15, 8, 36, -15, -46, 23, 31, -22, 39, -47, 24, 9, 5, -47, -32, 7, -1, -30, 38, -5, -17, 18, 36, 12, -12, 1, -34, -9, 27, 35, -10, -5, -41, 2, -21, 22, -12, -18, 13, 6, 38, -42, -39, -28, 8, -26, 43, -22, 33, -25, -5, -8, 5, 4, 40, 11, 35, -19, -6, -17, -21, 18, -25, 21, -28, -4, 35, 36, 4, -40, -13, 12, -28, -14, -41, 36, 17, 2, 42, -7, -15, -28, -32, -23, 1, -13, 29, -59, -44, -5, 45, -48, -19, -31, 19, -8, 28, 16, -33, 1, 36, -41, 0, 3, 45, -1, 4, 3, -5, -10, -5, -14, 27, 18, 15, -41, -3, 0, -1, 22, 28, 9, -45, 15, -8, 22, -13, -33, 11, 25, -8, 28, 43, 16, -26, -40, -18, -12, -19, -18, 39, -14, -17, 8, -32, -11, -7, 9, 15, 26, 19, -22, 48, -39, 42, 22, -28, 26, 23, -21, -39, 2, -2, -37, -2, 32, -32, -21, 44, -45, -21, -1, 35, -23, 20, 22, -14, 0, -15, -17, 6, 19, 3, -30, -25, -1, -8, -5, -36, -35, -21, 10, -3, -16, -21, -35, 6, -12, -15, 13, -9, 14, -27, -45, 33, -30, 35, -25, -27, 0, -35, 19, -36, -7),
    (12, -39, -48, 29, 59, 12, 14, 27, -42, 18, -14, 3, 18, -16, -22, 10, 5, 26, -54, 31, -35, -37, -10, -18, 13, 20, 23, 26, -16, -22, 50, 42, -6, -27, 14, -9, 10, -21, -7, 10, 2, -25, -17, -16, -5, -12, -44, 1, -17, 23, -9, -10, 5, -34, -43, -2, 47, 21, 1, 29, -32, -4, -25, 50, 33, -44, -20, 5, 12, -15, 25, -4, -38, 16, -24, -33, -6, -10, -28, 25, -22, -7, 7, -36, -10, 6, -34, 24, 6, 7, -9, 35, -14, -1, 33, -3, 3, 16, -20, 26, 51, 45, 15, -37, -39, 22, -17, -1, -39, 30, -13, -9, -34, 68, -17, 30, 13, 2, 1, 20, -8, 6, 22, -8, -44, 25, 3, -21, 17, -24, 12, -8, 30, -6, 20, -11, -54, 29, -55, 1, 32, -2, -43, 23, -37, 41, -33, 29, 29, -26, -7, -13, 23, 27, 43, 10, -45, -3, -5, 22, 25, -4, 32, 0, -4, -43, -6, 4, 4, -11, -14, 32, 41, 34, -18, -12, -1, 5, -39, -20, 8, 12, 3, -4, -33, 37, 23, 42, -14, -4, -7, -3, -26, 27, -4, 10, 44, -1, 17, -32, -9, 23, -9, -21, 1, -25, 17, -28, -10, 23, 28, -17, -3, 4, 19, -26, 4, 0, -20, -48, -20, 0, -21, -18, -33, -26, 4, -7, 27, 15, 11, -20, -3, 12, 7, 18, -20, 21, -11, -42, -22, 69, 13, 27, -16, -23, 46, -27, -23, 39, -10, -16, -19, 12, -6, -10, 29, -27, 1, -14, -13, -28, 5, -21, -3, 17, 25, -22, -31, 7, 19, -25, -29, 10, -41, -9, 19, -27, 23, -37, 28, 27, 5, 32, 9, 0, 20, -50, -3),
    (-5, 16, 7, -23, -27, 9, -23, 20, -17, -10, 17, -20, -52, -50, 36, -12, 6, 28, -8, 43, 16, 38, -37, -7, -46, 1, -77, -11, 15, -37, 9, -45, 16, -20, 21, 4, 15, -16, -14, -7, -39, -12, 20, -34, 5, -8, 21, -48, 10, 21, 40, -20, -1, 35, -17, -21, -53, -35, -17, -60, -30, -30, 2, -16, -7, 18, -16, -17, 38, 51, -9, 30, -7, -8, 24, -6, 2, -9, 13, -13, -22, 15, -6, -25, -50, -9, 23, -7, -34, 1, -11, 23, 56, -13, -28, 0, -6, -1, 30, 31, -37, 10, -25, 21, 10, 3, 44, -8, -25, 21, 19, 18, 14, 28, -30, -18, 25, 37, 16, 0, -29, -40, -46, -46, -28, -5, -16, -21, -21, -50, -13, 29, 23, -15, -51, 11, -5, 16, 17, 22, 0, -23, 3, -55, -17, 25, -1, 4, 1, 15, 40, -5, -26, -20, -42, -40, -20, -3, 12, 22, 6, -7, 23, 44, 12, 14, -11, -3, -3, 2, 5, -15, 24, 14, -22, -24, -24, 35, 26, 23, -23, -4, 41, 3, -22, 35, -35, 35, 35, 22, -20, -10, -3, -36, -10, -10, 1, 13, -52, 13, 12, -9, 13, -18, -34, -3, -2, -25, 20, 8, -4, -6, 37, 28, -11, -17, 36, -42, 3, -9, 22, -1, 7, 43, 19, -17, -25, 35, 43, 40, -5, 5, -7, -25, 65, 3, 3, 43, 16, -37, -8, 51, -27, -25, 4, -12, 48, -26, 32, -5, -64, -37, -3, 29, 49, 21, -14, -20, -25, -5, -8, -13, -8, 29, 26, -10, 36, 49, 21, 14, 3, -17, -27, 42, -33, 2, 45, 10, 19, -6, 32, 14, 12, 17, -15, 9, 21, -24, 39),
    (0, -20, -32, 7, 25, 12, 27, 15, -14, -22, 35, -23, -7, -2, -2, -33, -13, -2, -19, -38, 41, 28, 35, -14, -16, 17, -24, 4, -20, 22, 25, 1, 32, -30, -6, 40, 5, -4, 25, 20, -16, -9, 61, -11, -22, -11, -40, 16, 7, -9, -14, -40, 28, 45, 30, -12, 5, 30, -13, -23, -8, 19, -15, 39, -13, -4, 29, -8, -32, 16, 7, -13, 7, -14, 16, 4, -3, -16, -3, 16, -12, -5, -43, -12, 3, 29, 11, -28, 14, 38, -3, -47, -7, -32, 3, 31, 25, -65, -47, 20, 19, -33, 19, 1, -35, -56, 23, 7, -27, -9, 0, -21, 2, 3, -37, -26, 34, 24, 32, -35, -6, -12, -49, -32, -10, 13, -22, 63, 10, -34, 6, -21, -50, -5, 42, 40, -4, -5, 28, 0, -19, -1, -28, 6, 17, -27, -20, -46, 8, 2, -11, 6, -41, -14, -30, -24, -44, -25, 3, 10, -19, 18, 6, 37, -8, 20, 21, -1, -3, -9, 12, -45, -31, -17, 0, -58, -25, -50, -4, -22, 16, 56, -2, 34, -20, -1, -31, -50, -5, -7, -9, 3, 28, -26, -46, -6, 48, 15, 14, -20, -32, -11, 13, -6, 6, 19, 7, 37, -12, -35, -48, 11, -19, 11, 5, -19, -18, 6, -13, -12, 18, -37, -40, 29, -3, -54, 27, -2, -6, 31, 10, -13, -25, -7, 51, 5, -26, 13, -5, 4, 26, -17, -35, 10, 45, 18, -5, 29, -11, -3, -4, 22, 33, -26, 16, 27, -10, -19, -11, 49, 18, 12, 48, 45, 23, -39, -9, 16, -7, 17, 7, 8, -26, -28, -10, 19, -5, 12, -12, 43, -5, 43, 22, 1, 0, -5, -8, 38, 7),
    (-35, 38, -42, 22, 1, -6, 22, -20, -32, 28, -18, 18, 15, -16, -45, 38, -8, -17, 22, -11, -19, 3, -22, 11, 12, -15, -15, 18, 46, -3, -6, 3, -39, 17, -48, -33, -2, -51, 18, -11, -32, 13, 3, -14, -14, -24, 8, -6, -12, -56, -8, 23, 1, -4, 30, 9, 17, 22, -24, -13, 29, 20, -7, 10, 12, -10, 6, -25, 34, -4, -10, -9, 6, 31, -29, -30, -7, 31, 24, 24, -39, -37, -12, 26, 5, 4, 46, 15, -21, -21, -2, 40, -18, 24, -32, -18, 25, 20, 12, 14, -44, 3, 14, -1, 36, 51, 0, 33, 19, -15, 6, 16, 4, -23, -28, 10, -17, 5, -34, 1, 9, -34, -26, -13, 14, 21, 16, -6, -29, 25, -9, -21, 3, -7, 23, -26, 28, 45, -34, 21, 29, 14, 81, -22, -17, -24, 17, 50, -2, -17, 31, -8, -4, -5, -22, 7, 41, -23, -18, -21, 27, -25, 37, -5, -17, -36, -15, -19, 20, 9, -33, 8, -43, 27, 28, 15, 12, -14, 6, 11, -10, -27, 51, 2, -30, 40, 6, 19, 8, -47, -30, -19, 5, -9, -2, -31, -1, -37, -14, 6, -15, 17, 18, 2, 15, 2, 2, 22, -33, -60, 9, 3, -30, 13, -19, -19, -9, -31, 46, -15, 28, -46, -8, 18, 28, 23, 36, -27, -9, -16, -23, -5, 4, 30, -26, 32, 20, -41, 29, 22, -10, -11, -37, 30, 17, -31, 0, -27, -1, -12, -9, -21, 22, -24, -17, 13, -23, 2, 38, 28, -45, 11, 24, 19, 20, 36, -2, 4, 20, 1, 17, 19, -3, -20, 7, 2, -5, 23, -2, 28, 18, 16, -6, -10, 27, -11, 8, -18, 4),
    (-9, 43, 18, -35, 1, 19, 22, -3, -35, 19, -4, 50, 3, 30, -14, -5, 17, 10, 18, -20, -3, 1, 9, -43, -22, -7, 10, 19, 26, -24, 27, 37, 1, 21, -23, -40, -30, 14, 34, 0, 6, -21, -14, 25, 8, -16, -32, 9, 1, -4, 44, -39, 4, -26, -4, -37, 12, -21, 58, -24, -30, 15, 23, -23, -31, -6, -33, -33, 17, 33, -22, 1, -13, 8, -7, -4, 7, 21, -18, 2, 14, 19, 0, -13, 0, -18, -25, -42, -36, -32, -16, -31, -37, -30, -28, 28, -25, -1, 24, -38, -13, 24, -41, -8, -3, 20, -13, 8, -11, -22, 9, 41, 8, 0, -36, 3, 29, 45, 4, -51, 0, 32, -18, 53, -1, -41, -22, 2, -14, 12, 21, -4, -40, 18, -7, -12, 20, -27, -40, 28, -39, 16, 25, -9, -14, 18, 30, -15, -15, 49, -29, -52, -12, 0, 14, 17, -8, 21, 28, 36, 8, -9, 18, -33, 6, 28, 0, -2, -37, 6, 15, 18, -41, -18, 23, -20, -11, 3, -20, -60, 7, 24, -21, -30, -34, 11, -5, -18, -3, -37, -36, 23, 15, -4, 33, -12, -4, -15, 5, 21, 26, 32, -46, -20, 12, 4, 2, 12, 5, 10, 25, 30, -6, 5, -38, 5, -39, 7, 5, 47, -3, -18, -2, -4, 47, 11, -11, 15, 5, -7, -14, 9, -2, -15, -68, 5, -22, 10, -2, 44, -18, -44, -7, 2, -12, 59, -6, 8, -10, 12, -30, 7, -4, -18, -20, 23, -11, 8, -25, 1, 31, 24, 6, -37, -28, -22, -11, 35, -63, -11, -2, 0, -21, -58, -47, -33, -15, 38, 36, -31, 17, -6, -4, -35, -4, -31, -6, 17, 3),
    (-26, 26, 41, -7, -11, 30, 11, -29, -5, 4, -61, -22, -20, -21, -30, -7, 1, -10, 23, -43, -6, 11, -24, -11, 19, 8, -19, -22, 9, -2, -5, -14, -2, 30, 60, 25, -37, -25, -6, -69, -35, -20, -49, -26, 4, -2, 11, 20, -33, -37, 16, -23, -43, 55, 14, 27, 40, -23, 40, -22, -18, -11, 52, -26, 14, 12, 31, 24, 13, -25, 2, -39, 16, 11, -17, -16, -37, 8, -19, -27, 11, -13, -9, 11, -15, 1, -24, -16, 40, -59, 46, -18, -3, -4, 53, -21, 23, 28, 24, 3, -32, -4, -29, -39, 12, 15, -34, -13, 20, -34, -24, 17, -6, -42, 23, 12, -35, 5, -7, -57, 40, 0, 52, -51, -12, 20, -35, -53, 23, 2, 18, -25, -42, -11, -29, -30, 2, -10, -8, -35, -36, -34, -30, 34, -44, -71, 25, -7, 6, 33, -23, -6, 16, -49, 20, -5, 41, -30, -35, 26, 21, -49, -39, -8, -16, -33, 2, 2, -20, -16, 36, -22, -57, -33, 36, 6, -6, -58, 28, -28, -22, -26, -21, 19, -11, -51, -8, 42, -20, -16, 26, 46, 10, 4, -25, -20, -12, -34, -11, -11, -24, 8, 13, 26, -7, 12, 22, 32, 11, 17, 7, -15, 31, 11, 29, -6, 7, -37, -25, -21, 14, 33, -10, 14, 23, 2, -10, -18, -10, -42, 0, -21, -36, 8, 3, -42, 8, -20, 12, 4, -31, -1, -34, 16, -20, 18, -25, -32, 28, 30, 10, -10, 12, 31, -16, 16, -11, -9, 17, 0, -1, -14, 9, 20, 6, -31, -15, -34, -5, 6, 36, -54, -14, -15, -21, -41, -10, 13, -48, -17, 5, -4, 5, -5, 35, 15, -32, -33, -5),
    (-26, -23, -28, 9, 11, 41, -51, 14, -20, 4, 2, 23, 40, -29, -36, 40, 10, 2, -56, 15, 9, -71, -29, -11, -48, 19, 25, 13, -25, -21, 33, -15, 7, -25, 11, -11, 13, 27, 13, -19, -19, 1, -15, -26, -11, 4, 13, 36, 44, -8, 3, -21, -3, -15, -25, -7, -30, -19, 47, 25, 10, 0, -7, 3, -19, -33, -3, 8, -13, 10, 7, 27, -39, -19, -52, 22, 24, 37, 20, 11, 35, -23, -2, -25, 12, 17, 12, 16, 2, -7, -18, -45, -9, 8, 25, 8, -2, -2, 36, -23, 13, 7, -39, -10, 24, 14, 0, -43, 3, -16, 25, 48, 27, 14, -5, 41, -30, -14, 2, 12, -45, 30, -30, 16, 34, 3, 33, -30, 28, 15, 60, -11, -21, -47, 7, -21, 19, 21, -64, -18, -26, 26, 31, 26, 4, 8, 44, -14, -14, -19, 19, 28, -10, 13, -10, 12, -6, 23, 3, -58, 5, 34, -7, -29, -8, -20, 23, -44, -5, 38, -31, 20, -23, -16, -15, 47, 11, 8, 31, -21, -4, 5, 3, -24, -10, -17, 16, -38, 12, -25, 5, -61, -18, -6, 33, 0, -30, -20, -9, 27, 27, 9, -19, 10, -17, -12, 5, 23, 4, 22, -8, 14, 12, -6, 14, -14, -4, -27, -49, 9, -35, -8, -22, -50, -25, 37, 26, 4, -7, -4, -41, -22, 6, 24, -39, -3, -37, -47, 11, 12, -3, 11, 35, 19, -36, 6, 13, 26, 8, 9, -19, 9, -29, 21, 25, -75, -20, 26, -39, 19, 20, -29, -25, -3, -20, 11, 19, 23, -40, -13, 16, 26, 24, 9, -27, -32, -3, 14, -7, 24, -32, 12, 10, -7, -8, -14, -32, -24, -3),
    (23, -1, -2, 7, -16, -62, -39, 25, 14, -10, -22, -1, -30, 2, -2, 29, 55, -35, 42, -35, 3, -16, -48, -24, -10, 5, -20, -16, -26, -24, 1, -27, -1, 1, 34, 8, -13, -31, -46, -25, 3, 1, -5, -19, -3, 27, 56, -21, 33, -23, 17, -61, -15, 4, 16, -23, 21, -20, -20, 0, 1, -12, -13, -40, 16, 0, -1, 15, -12, -25, -19, -49, -39, 20, -5, 12, 1, 25, 25, 23, -37, -27, -37, -31, -31, 12, 13, 22, -8, -3, -36, -20, 36, 12, -15, -8, -9, 21, -8, 22, -18, -26, -45, -25, -9, -39, -13, -12, -33, -11, 21, -37, 26, -13, 36, -24, 5, -5, -22, 9, -53, -19, -36, -7, -21, -28, 21, -34, 12, 13, 41, -18, -12, -7, -62, 10, -60, -32, 31, -31, 5, 30, 71, -11, 57, -8, 5, -27, 9, 11, -29, -16, -8, -36, -30, -37, -12, -36, 17, -29, -20, 3, 21, 8, -10, -34, -35, 14, -24, -15, 28, 22, -31, 34, 74, -29, 27, 7, -3, -58, 25, 44, -6, 24, -21, -6, -53, -11, 13, -24, -1, -23, -9, 57, 6, -21, -19, 24, -16, -32, -4, 12, -14, 22, 9, 0, 21, 42, 13, 23, 27, 2, 38, -15, 33, 22, 8, 26, -1, -18, 11, 1, -6, -4, 10, 57, -6, -15, 17, -28, -37, -26, -46, -8, 4, -45, -8, 17, 29, -14, 32, 12, 30, 32, 34, 19, 10, 11, -18, -24, -26, 3, -38, 7, 0, -6, -8, 0, 16, 13, 38, -34, -32, -5, 14, 0, 30, -33, 19, -17, 28, -23, 22, 21, 11, 13, -9, 8, 18, 25, -5, 7, -15, 12, -26, -53, 27, -25, -1),
    (19, -12, -27, -5, 16, 11, 15, 49, -6, 12, -48, 14, -21, 9, -28, -2, 27, -34, -3, 14, 4, 5, -1, 20, 8, 18, 13, 11, 37, 46, -17, 24, -1, 6, 36, 5, 36, -44, -4, 30, 16, 45, -54, 31, 6, 50, -53, 25, -4, -16, 25, 0, 24, 36, 32, -2, -26, 11, -8, 17, -4, 42, -26, -56, 29, -28, 23, 7, 0, -43, 18, -17, -23, 13, -32, 24, -7, 26, -6, 30, 3, 5, 19, 29, 23, 54, 38, -8, -25, 39, 13, -11, -1, 11, 35, -35, -15, -36, 2, 4, -29, -13, 8, -24, -2, 14, -47, 29, -15, 21, 13, 35, 8, -61, 0, -20, -30, 9, 8, 21, -49, 23, -17, -24, 30, -20, -4, 19, -19, -13, -18, -11, -29, -32, -18, -37, -39, 17, -16, 6, -51, 8, 39, 13, -24, -36, -10, -32, 34, 41, 31, 18, -7, 31, -55, -60, 29, 3, -46, -16, 13, -20, 34, 18, -7, -44, -7, 4, -9, -48, -29, 18, -30, -46, 20, 24, -20, -17, -7, -23, 1, 15, -11, 6, 6, 25, -38, -8, -6, -4, -33, -34, -10, -61, 12, 21, -10, 3, 18, -29, -14, 18, -12, 12, -44, 7, -13, 39, -24, 21, 6, 13, 16, -57, 2, 21, -11, 1, -50, 1, 24, -34, -30, 31, 2, -8, 5, 47, -22, -23, -9, -29, 11, -19, 4, 5, -5, -41, -6, -1, 25, -37, 24, -22, -23, -13, -13, 50, -9, 21, -43, -29, -4, -26, 3, -7, 7, -34, 13, 37, 55, 12, -27, 18, 24, -30, 26, 1, 4, -25, -7, -4, 11, 8, 2, -23, 15, 7, -9, 24, 12, -18, -59, -16, 18, 40, 27, 30, 0),
    (-7, -2, 3, -20, -31, 6, 16, -19, 20, -15, -45, 28, -33, -11, -6, 16, -18, 25, 2, 16, 4, -1, -7, 6, 31, 40, -32, -16, -8, -6, -1, 5, -11, 11, -3, -10, -30, -21, -29, -16, -10, 19, -16, -26, 15, -20, 42, 14, -29, 70, -35, 30, 16, 25, -21, 19, 29, 34, -32, -29, -12, -45, 27, -1, -12, 3, -2, -16, -5, -38, 21, -16, 15, -13, -2, 13, -43, 8, 48, -1, -38, 48, -41, 40, 11, 16, -22, 31, 54, 36, -32, 1, -17, 25, -22, 9, -40, 0, -19, 11, -17, -26, 6, -12, 17, 13, -8, -33, -60, -1, 38, 37, -9, 64, -22, -14, -15, -3, -35, 40, 30, -37, 3, -2, -26, -13, 4, 25, -11, -8, -18, 0, -28, 6, 19, 30, 26, -31, 52, -22, -36, -28, 31, 23, -27, 102, -24, 22, -16, 3, -15, 27, 25, -20, -7, -3, -43, -21, 8, 11, -24, -4, -39, 3, -8, 10, -14, 27, 44, -46, 46, -42, 13, -10, 28, -20, 5, 44, -14, 27, 13, 19, -33, 11, 14, -8, 7, 52, -37, 19, -49, 0, -31, -26, -19, -9, -9, -37, -17, 45, 2, -25, 6, -38, -1, -46, 3, 10, 9, 5, 25, 28, -15, 12, 2, 40, -24, -40, -14, 44, -8, -22, 7, 10, -20, -23, 3, -10, 10, -23, 8, 22, 8, -17, 15, -25, -16, 9, 30, -2, 23, 29, 5, 53, -2, -42, -7, 48, 5, -3, -13, 7, -56, 17, 6, 5, -33, 6, 4, -29, 12, -23, 10, -42, -19, -51, 10, -46, 32, 4, 12, -15, 2, 41, 12, 7, -4, 13, 17, -3, 2, 15, 14, 2, -11, -11, -7, 14, -6),
    (-9, 6, -20, -26, 20, -7, 22, -40, 17, 35, -33, 2, 31, -23, 3, 18, 13, 30, -14, 4, 40, 39, 21, -7, 2, -11, -23, -21, -67, -23, 35, -41, -27, -16, 30, 8, -9, -19, 25, -32, 0, -16, -37, -11, -15, 12, 33, -17, 4, 59, -13, -25, 17, 14, -15, 4, 31, -51, 21, -58, -29, -32, 36, -7, 20, 28, 24, -7, -8, -17, -3, -33, -3, 33, -57, 10, -1, 17, 13, 42, -15, 36, 6, -63, -20, -15, -13, -23, -1, -50, 17, -24, -45, -2, 27, -37, -11, 30, 27, -44, -3, -3, 51, -37, -26, 5, -25, 6, -15, -29, 14, -16, -9, 23, 40, -3, -28, -22, 14, 21, -14, -62, -15, 22, -44, -44, 34, -36, -13, 51, -4, -11, 0, 10, 10, -7, 14, 33, -27, -29, -17, 20, 11, 30, -8, 35, 40, -58, -26, 1, -19, 7, 16, -19, 36, -3, -19, -24, 37, 6, 17, -2, -5, -20, -7, -21, 46, -28, -8, 31, -36, -1, -1, 28, 21, 31, 24, 2, 36, -61, -19, 31, -20, 23, 13, -37, 23, 35, 8, -2, -2, -10, 27, 8, -3, 8, -10, 7, -23, -39, -20, 26, -3, -16, 41, 21, 7, 28, 26, -2, -5, -36, -33, -25, -11, 10, 0, -17, -4, 22, 39, -8, -4, -31, -21, -17, 10, 20, -32, 35, -61, -12, -5, 38, -22, 17, -9, 8, -37, -1, -1, -69, 32, -39, -2, 6, -51, -23, 2, -2, 35, 1, 25, -60, -24, -36, 5, -32, -8, 5, 35, 46, -6, -12, 1, 6, 4, -27, -14, 10, 23, -25, 12, -68, 44, -32, -15, -26, -40, -9, 30, -13, -19, -5, 35, 2, -72, -23, -2),
    (-15, 17, 14, 22, 14, -3, -16, -15, 2, 38, -22, -35, -43, 59, -23, 30, -29, 35, -10, 5, 10, -14, 5, 27, -17, -12, 33, -4, -5, 10, 45, 35, -6, 6, -15, 6, -6, -9, 0, -19, 18, 48, -9, -38, -21, 73, -50, 21, 13, 50, -48, 15, -5, -11, -11, 24, -2, 3, 13, 11, 30, 53, 30, 19, -9, 18, 19, 13, -16, 0, 19, 14, -13, 54, -25, 11, -1, 35, -59, 27, -28, 18, -31, -5, -15, -16, -20, 38, 1, 32, 27, 33, -3, 21, -8, 21, 5, -35, 18, 8, -42, -25, 9, -35, -24, -20, 8, -35, -6, 20, 27, -6, 17, -9, -35, 5, 29, -1, 4, -16, -6, 21, 12, -26, -32, -20, 26, 1, -26, 26, -18, 14, -12, 13, -27, -24, -4, 23, 69, -32, -10, 30, 16, 5, -47, 15, -30, 14, -24, -14, -5, -13, -12, 30, -11, 17, 18, 26, 46, 28, -17, 12, -9, -20, -31, 31, 8, 12, 3, 30, 0, 6, 23, 45, -21, -19, -43, 33, -44, 10, -36, 2, 12, 28, -2, -15, -32, -16, -19, 28, 18, 6, 5, 17, -19, -38, -33, -17, -34, -4, 23, -7, 8, -30, -1, 35, 21, -29, 16, -15, 20, -1, 19, -52, -50, 23, 24, -41, -20, 45, 10, -49, -4, 27, -17, 21, 25, -26, -35, -5, -11, -8, -10, -33, 46, -28, 18, 36, 36, -42, 9, -39, 19, -10, -38, -12, -42, 4, 32, 4, -38, 26, 13, -62, -21, 42, 3, 31, -9, -16, 13, 5, -10, 13, 15, -5, 25, -14, -25, -22, 12, -12, 9, 32, -42, 25, -29, -5, -26, 10, 21, -22, -39, 1, -9, -26, -12, 32, -10),
    (25, -17, -15, 30, -3, -6, 24, 10, -4, 19, 7, -11, -25, 31, 20, -31, -32, 24, -12, 1, 32, -19, -10, 9, -2, -2, -33, -50, 24, 37, -2, 10, -5, -35, -34, -9, 25, 37, -27, 3, -8, -1, -33, -6, -9, 25, -20, -18, -12, 47, -11, 2, -26, -19, 25, 29, 40, -54, 2, 1, 23, 20, -7, 57, 5, 8, -29, 7, 28, 1, -22, 25, 48, 14, 12, -34, -2, 11, -3, 6, 33, 27, -22, -36, -25, -50, 18, 32, 22, -13, 26, 34, 1, 14, -7, 65, -27, 4, -27, 14, 26, 62, 20, 31, 37, -27, 30, 10, -36, 12, -35, 9, -18, 18, -9, -45, -50, -45, -2, -19, 37, -31, -45, -30, 49, 28, -14, 49, -13, -13, 23, 17, 25, 24, 14, -8, 11, -44, 9, -41, -20, 45, -14, -18, -3, 16, -30, -9, -19, -48, 3, -9, -24, -7, 35, -22, 16, -1, 17, 45, -54, 11, 29, -13, 24, -14, 27, 5, 25, -10, -1, 8, 5, 7, 9, -34, 6, -1, 17, 9, 1, -43, -8, 35, 1, -20, -2, 13, -36, -20, 4, 17, -24, -21, 7, -28, 3, 4, 26, -4, 51, -25, 28, -10, -1, -24, -6, -38, -27, -18, -4, -47, -16, 34, -22, -20, -2, 17, -54, 0, -39, -28, -34, 19, -11, 25, -22, -39, -50, -3, -6, 27, 18, -34, 6, 21, 7, 0, -8, -35, 4, -51, 2, -9, -6, 9, -24, -45, -27, 5, 12, 35, -18, -10, 12, 3, -4, -8, -44, -20, -35, -23, -12, 27, -30, -41, -9, 24, -1, 32, 15, -2, -20, -9, 33, 7, -11, 11, -10, 3, -39, 20, -25, 23, -28, -29, -29, -22, -7),
    (9, -16, -16, -22, 22, 28, -31, -36, -4, -25, -13, 8, 22, -23, 8, 33, 36, -21, -9, 14, 31, 31, -6, 12, 28, 27, 17, -10, 3, 30, 3, 26, 32, 12, -24, 17, 40, 24, -36, 1, -35, 27, -12, 13, -25, -14, -14, 5, 12, -5, -2, -14, -3, 40, 8, 19, 18, 50, 1, -16, 20, 13, 17, 25, -20, -16, -34, -14, 23, 8, -1, -11, -1, 7, 15, -7, 24, 11, -12, 21, 3, -16, 0, 11, 23, 45, 15, -17, 28, 4, -21, 14, -20, 45, 24, 8, 35, -34, -14, 3, -1, 17, 22, -47, -18, 22, -5, 27, -21, 20, -34, 1, -31, -42, -4, -26, -4, -24, 6, 23, 29, 21, 19, -8, 19, 59, -20, 3, 24, -43, -25, 44, 16, 50, -19, -12, -46, 15, -46, 55, 5, 18, -40, 42, -31, -44, 4, 20, 16, 30, 21, 3, 12, 8, 23, 13, 13, 34, 6, 18, 21, -40, -20, 14, 44, 10, -12, 14, -6, 26, -29, 18, -26, 50, -15, 30, -22, 0, 1, 6, 9, 46, 1, 3, 30, 2, -2, 53, -26, 29, 27, -14, -35, -65, -13, 26, 13, 35, -44, -31, -38, 1, 33, 24, -19, 43, 22, -31, -25, -37, 19, 12, 8, 16, 40, -43, -17, -11, -4, -61, -11, 19, 17, 26, 11, -39, -20, 10, 30, -30, -21, -48, 8, -22, 18, 28, -1, -13, 28, 38, -31, -29, -2, -7, -9, 7, 18, -11, -12, -26, -21, 19, 17, -9, 13, 14, 1, -4, -20, -6, 53, -47, -19, 13, -28, 16, -2, 0, 12, 18, 7, 1, -25, 11, -9, -34, -33, -11, 23, 31, 6, -6, -6, 2, -25, -7, 17, 1, -8),
    (3, 33, -19, -12, 18, 31, -28, -41, 7, 26, -50, -33, 7, 5, 18, 2, 49, -32, 29, 47, 22, -22, -18, -24, -32, -30, 11, 47, 22, -40, 8, -7, -19, 3, 39, 24, -20, -9, -61, -26, -12, 20, -18, 14, 9, -37, 33, -28, 17, -25, 4, -34, -21, -41, -13, 24, -47, 16, -5, -3, -6, -50, -12, 32, -2, -9, -17, 3, -20, 17, -40, -2, 14, -28, -26, -40, 3, 0, 20, -34, 13, 13, 31, 3, 24, -24, -25, 16, -23, -36, 4, 16, 14, 19, 11, -19, -20, 10, 17, 9, -33, 57, -36, -3, -36, 15, -10, -4, 21, 28, -33, 6, 24, -7, -12, -2, 11, -55, 21, 0, -18, -33, 20, 21, -23, 29, 28, -28, 38, -17, 40, -43, -55, -2, -16, -31, 14, -23, -59, -2, 19, -13, -13, 29, -12, -32, -1, -32, 29, 3, -6, -3, -61, 18, -30, 26, 16, -36, -17, -45, -8, 40, 43, -22, -33, 3, -28, -25, -27, 33, -30, -27, -20, 36, -1, -20, -5, -18, -6, 2, 14, -47, 9, 11, 18, 1, -24, -20, 3, 1, 35, -27, 3, 42, -33, 5, 22, -8, 11, 9, -12, -13, 5, -10, -4, 6, 9, 30, 15, 2, -13, 47, 24, 2, -21, -34, -22, 0, -10, -22, 24, -33, -3, 33, -28, -2, 19, -43, -23, 23, -25, -18, -31, -22, -5, -26, -36, 37, 20, 19, 31, 27, -29, -8, -18, -42, -13, 33, -47, -25, -20, 23, -42, -31, 28, -20, 11, 40, 45, -52, 10, -1, -18, 1, -40, 30, -24, 12, 11, -2, -12, 8, 25, 13, 14, 8, 23, -57, 21, -23, -33, -29, -12, 27, 3, -5, 17, 6, -1),
    (-31, -20, 13, 14, -36, -10, -14, -24, -3, -39, 60, -34, 12, 6, 37, -9, 26, 25, -24, -51, -6, -44, 2, -31, -6, 6, -26, -39, -27, -63, -22, 39, -43, -42, 17, 3, 32, -10, 3, -39, -4, -18, 37, -42, -9, -23, 60, -32, 18, 30, -23, 16, 22, 0, -25, -35, 22, 4, -2, -34, 24, -26, 3, -6, 7, -30, 41, -9, 7, 5, 2, -50, 12, 14, 34, 25, -3, -33, -2, -4, 43, 38, 10, -7, 22, -22, 18, -34, -10, -22, -18, -51, 5, 16, 20, -25, -50, 29, 4, -4, -25, 5, -28, 29, -23, 36, 13, 10, 45, -19, 9, -45, 7, 19, -27, -7, -35, -4, -16, -35, -48, -30, 42, -31, 14, 18, -25, 22, -36, 34, 33, -2, 14, 1, 30, 37, 28, -11, 56, -18, 39, -11, 0, -30, 20, 62, -1, 26, 25, -19, -2, -18, -20, -11, 23, -15, 12, -15, 35, 41, 4, 4, 18, -30, 35, 3, 17, 15, -11, -15, -7, 32, 25, -4, 13, -11, -14, 26, -35, 37, 25, -24, -4, 11, 17, -25, 36, 5, 12, -2, 23, 40, 20, -2, -17, 6, -4, -8, -8, 14, 4, -23, -29, -32, 37, -14, -32, 7, -19, 13, 16, 20, -12, 3, 18, 2, -22, -12, 23, 29, 9, -33, -7, 40, -3, -11, -17, 39, 16, -12, -17, 31, -19, 22, -13, -8, 2, 36, 2, -2, 5, -10, -16, -23, -30, 10, 15, 1, -45, 4, 21, 21, 9, 26, 35, 59, 12, 9, -30, -13, -20, -2, -20, 30, 2, 29, 6, 26, -10, 11, -2, 0, -4, 11, -30, 6, 28, 28, -18, 17, -36, -40, 12, 10, -27, -5, 30, 13, 9),
    (-24, 36, 31, -10, -54, 35, -11, -16, -31, 7, 18, -50, 3, 11, 22, -26, 21, -8, -28, 17, -4, -12, 11, -24, -17, 23, -36, -20, -4, 16, -23, -25, 16, 24, 20, -7, -2, 43, -21, -29, -19, 25, -4, -12, -26, -28, -27, -27, -39, 0, 5, -5, 11, -5, 24, -15, -6, -3, -27, 12, -14, -16, 62, -33, 15, 10, 2, -15, -21, 27, -8, -15, -41, 34, -45, 2, 14, 7, -3, -15, 38, 23, 14, 20, 30, -46, 0, 8, -2, -19, -1, 4, -4, -5, 31, -41, -49, 8, -9, 0, -26, 35, -71, 31, -17, -2, 43, -43, 16, -32, 24, -19, -18, -22, 37, 0, 8, 14, -1, 24, -34, -6, -10, -3, -34, -17, -2, 26, -23, 45, 11, 10, 2, 37, -37, 12, -2, 16, 24, -32, 38, -34, 39, -11, 13, 31, -34, 6, 6, -41, -17, 17, 1, 23, 0, -25, -12, 1, 39, 31, -24, 58, 27, -44, -16, 19, 6, -8, -21, -8, 10, 29, 41, -2, 30, -2, -8, 51, -33, 1, -6, -44, 11, -22, 17, 13, -7, 14, -8, 21, 44, -2, 24, -36, -40, -9, 23, 12, 37, 10, -1, 21, -42, -2, -28, 24, -20, 8, 25, -15, 29, 11, 4, -1, 5, -8, 4, 19, -29, -8, -27, 5, -29, -10, 1, -28, 3, 23, 3, -1, 17, 18, 35, 44, 19, -6, 44, -35, -5, -19, -21, -24, 22, 23, -3, -5, -17, -19, -27, 34, -10, -19, 14, 24, 6, -8, 13, 17, 3, -27, 7, 40, 36, 20, 21, 29, -28, -27, 31, -25, 10, 29, -31, 15, -7, -24, -48, -9, -5, -5, -21, -4, -9, 21, -26, -24, 0, 3, -2),
    (9, 23, -13, 14, -21, 5, -17, 17, 11, -16, 11, -25, 39, -8, 31, -29, 21, -19, 28, 24, 26, 10, -13, -2, 14, -10, -15, 17, 23, 32, -43, -17, -47, 45, 10, 4, -22, 9, 14, 12, 15, 40, 22, 10, 33, 38, -30, 16, -10, 25, 4, -14, -27, -18, -15, -19, -8, 18, 0, -30, 9, 19, 18, -2, -34, -12, -24, -16, 5, 17, -13, -9, -22, 29, 17, 9, 29, 31, -25, -11, -11, -30, 5, 4, 13, -36, -25, -30, -10, -29, 1, 0, 43, -16, 29, -10, -20, 0, 27, 32, 33, 14, 41, 31, -5, 17, -5, 6, 35, 4, -41, 22, -4, -46, -13, 13, -1, 23, 19, -23, -20, 20, 72, 27, 5, 42, -27, 7, 39, 49, -45, -1, 17, 34, 24, -22, -18, 3, -35, 20, 32, 20, -48, 18, -13, -35, 3, -20, 25, 2, 15, -2, -56, 10, 8, 24, 27, 43, 21, 48, 28, -24, -15, -30, 11, 12, 6, 5, -1, -11, -4, -4, -5, 8, -27, 19, -4, -10, 11, -12, -12, 3, -8, 3, -58, 29, -7, -42, 7, 26, 36, 2, -12, -4, 12, 45, -12, 39, -18, 36, -2, 13, 16, 1, -6, -29, -37, -21, -22, 1, -31, 45, 5, 3, -13, 13, 10, 40, 8, 6, 2, 3, -26, -14, 24, 32, -5, 12, -12, 22, 15, -16, -28, -26, -6, -8, 34, -28, -25, -28, -35, -38, -13, 1, -9, 46, 35, 9, -10, 38, -39, 34, 32, -2, -26, 1, 22, 6, -35, 30, 17, -39, 9, 26, 15, -34, -41, 0, -19, -6, -18, -1, -1, -41, -35, -39, 17, 70, 34, -6, -24, 40, -19, 23, -5, -25, -30, -17, -1),
    (2, 23, -4, -13, 38, 34, -11, 0, -9, -26, -20, 29, 19, 14, 0, -15, -45, 14, 5, 5, 14, -51, 18, 4, -26, 57, -3, 44, -25, 38, 17, -25, 46, 21, -10, -1, 24, 17, 21, 14, -2, -18, -17, 44, 34, -28, -32, 34, -59, -1, -26, 0, -15, 1, 17, -9, 16, 40, 23, 42, -19, 24, 7, -43, 33, 21, 25, -22, 14, 31, 4, -27, -2, 0, -7, 37, 28, 17, -34, 1, -30, -25, -1, -29, 11, 5, 23, 25, -22, 50, 36, -8, 27, 21, 5, -25, -8, 21, 16, -22, -36, -35, -56, -28, -5, 6, -21, 0, -11, -12, 23, -12, -19, 45, 13, 9, 0, -28, 15, -18, 1, 50, -41, 40, 28, 19, -20, -50, 60, 8, 29, 6, 3, -26, -18, 3, -52, -25, -11, 4, 18, -13, 1, 2, -18, 13, -2, -22, -1, 33, 12, -34, 1, 78, 5, 9, -9, 17, 7, -13, 46, -19, 16, 21, 7, -3, -2, 3, 13, 16, 13, 30, 10, 11, 9, 6, -30, 8, -17, 24, 29, -9, 28, 2, -14, 16, -57, -27, 28, -2, -21, -3, 30, -35, 8, 11, -24, -6, -42, -16, -35, -39, -5, -4, 3, -56, 9, 3, 24, 51, -19, 11, 18, -13, -18, 0, -29, 13, -8, -26, -31, -27, -10, -20, 13, -6, -28, 25, -44, -70, -41, -25, -38, -19, 37, 7, -33, 4, 20, -4, -55, 36, -71, -5, 26, 41, 23, 48, 20, 25, -6, -31, -39, 18, -4, -15, -26, -5, -21, 32, 8, -52, -30, -40, 1, -46, 36, -3, -5, -21, 20, -20, -32, 40, -65, -19, 20, 16, 22, -21, 8, -39, -20, -18, -45, -15, 7, -15, -3),
    (7, -11, -19, -31, 21, -1, -3, 23, -47, 33, -38, 7, 15, -6, 10, 16, 18, -7, 37, 34, 0, 1, -42, -14, -22, -18, 0, -6, -9, 4, 22, -3, 11, 27, -9, -9, -2, -1, -17, -18, 18, 15, -42, -10, -31, 42, -1, 35, 5, -24, 22, 3, 1, 2, -26, 25, 6, -10, 24, 31, -28, 6, -22, -54, -22, 27, 31, -35, -27, -14, -15, -25, -11, 19, -27, -17, -14, 29, -5, 47, -20, -4, 1, 0, -22, 22, 30, 11, 36, -12, -20, 36, 37, 6, -3, -40, -5, 18, 13, -39, 20, 15, -44, 4, 6, -27, -50, 32, -13, 17, -6, 44, 17, -16, 13, -5, -17, -52, -48, -1, -18, -6, -5, -3, 4, 10, 9, -24, 38, 47, 7, -19, 0, 6, -46, -17, -30, -11, -46, 15, 7, 36, 11, 36, 34, -67, 19, -37, 29, 20, 14, 6, -6, -32, 6, -31, 6, -4, 28, -56, -18, 3, -20, -6, -40, -46, -51, -33, -21, 56, -18, -52, -13, -20, 2, 16, 1, -36, 19, -16, 20, -1, -4, -31, 28, -7, 6, -31, 9, 25, 17, -39, 8, -22, -40, -23, 14, 28, -36, 25, -35, 20, -25, -4, -4, 14, 2, 3, 37, 10, -1, 30, 30, -23, -43, -15, -18, -20, 40, 27, 8, 27, -30, 15, -15, 23, 15, -9, -7, 13, -17, -20, -32, -21, 4, 2, -6, 14, -8, 31, -7, -26, 17, -19, 15, 37, 23, 1, -21, 19, -35, 8, -14, 44, 3, -7, 4, 5, 31, 15, -34, 16, 12, 3, 4, -11, -32, 25, -20, -14, -20, 13, -42, -40, -2, -19, 14, 41, -39, 30, -15, 9, -54, 23, -9, 18, 31, 22, -3),
    (-25, -21, 2, -24, 41, -18, -47, 38, -36, 13, 22, -6, 1, 28, 8, -8, -27, 14, -59, 6, -38, 20, -10, -17, -52, -16, -22, 34, -29, -66, -68, -19, -46, -19, -26, -40, 8, -9, -41, -14, -48, -43, 38, -15, 7, 1, 26, -8, 2, 22, -4, 47, -43, 33, 20, -28, -1, 18, -10, -13, 14, 3, -6, -4, -21, -46, 23, -10, -17, 6, 5, 24, 8, 9, 13, 24, -26, -26, 44, 19, 11, 28, -9, -8, 4, -16, -31, 31, -24, -23, 19, -5, 0, -23, -16, -8, -5, 51, -3, 33, -4, 24, -51, -15, -5, 29, -18, -28, 25, 6, 24, -28, -2, -14, -26, -25, -25, -14, 43, -19, 25, 37, 10, 37, -15, -24, -27, 2, 3, 8, 31, -1, 37, -19, -32, 6, -7, -28, -1, 4, -20, -30, -10, -20, 20, 12, 7, -41, 31, -31, 27, 31, -37, 2, -18, -13, 22, 15, -30, -46, -22, -4, -4, -7, 3, -16, -11, -3, -35, 11, -38, 14, 0, 20, 5, 11, 6, -11, -14, -4, -4, -1, -2, 11, -42, 27, 18, -48, -16, 8, -24, -44, 35, 23, 9, 2, -25, -45, -1, -1, 31, 15, -19, -15, -4, -27, -12, -11, -6, 32, 2, -24, 32, -11, 41, 30, 8, 0, -8, -20, -14, -25, 36, 3, 11, 6, -11, 35, -9, -64, -46, -16, 5, 17, 8, 26, -13, 0, 0, 1, 32, -68, 57, 15, -6, 8, -7, 32, 6, -10, -14, 17, 21, 15, -14, -40, 32, -47, 18, -17, 41, -69, -55, -26, 20, -20, 32, -10, -40, 16, -12, 3, -20, -62, -6, -30, -25, -29, 14, 24, 8, 19, -38, -26, -29, -23, -3, -39, 6),
    (-24, -55, -5, 15, 32, -30, 4, 4, -2, -18, -42, -2, 23, 37, -18, 30, -25, 33, -38, 24, 13, 9, -42, -5, 40, 9, 6, 38, -6, -1, -24, 0, 26, -54, -10, -39, -18, 1, 44, 27, 21, -29, -35, 12, 65, -6, -53, -8, -29, -4, -50, -8, 9, 36, -5, -7, -23, 21, 51, 31, -4, 5, -7, 21, 7, 10, -4, 20, -14, 27, 36, 1, 38, -13, -41, 37, 30, 14, -9, 14, 0, -29, -17, 16, -10, 1, 1, -4, -6, 19, 32, -40, -5, 16, -8, -10, 20, -16, 13, -28, 10, 18, 5, 19, -27, -12, -44, 6, 7, 26, -5, 2, -23, 2, -29, -8, 1, 5, -28, -18, 35, 33, 24, 54, -41, -21, -9, -40, 27, -24, -31, -18, 3, 15, 37, -3, -3, -5, -69, 5, -10, 47, 10, 1, -10, 37, -61, 51, -2, 0, -24, 16, 9, 7, 40, 64, -26, -17, -7, -4, 4, -45, 37, 19, -26, 21, 33, 15, 33, -3, -7, -17, 35, 1, -23, 21, -43, -20, -10, 24, -32, 37, -8, 26, 25, 46, 47, 49, -12, -1, -19, 13, 1, -5, -1, -38, -40, 37, -25, -27, 14, 15, -50, -9, -14, -1, -22, 19, -30, 29, 18, -15, 13, -7, -21, 2, 14, 11, 30, 25, 1, -11, 15, -9, 9, 17, -24, -5, 27, 18, -25, -28, -26, -42, 20, -24, 4, 21, 20, 36, -41, 30, -20, 44, -7, -25, -33, 18, 25, 22, 24, 12, 1, -7, -18, -21, -11, -17, -29, -11, 10, 28, 8, 15, -10, 11, -50, -12, 16, -19, -9, 19, -35, 19, -39, -12, 6, 22, -4, 5, 3, 24, 12, 20, -55, -12, -1, 25, -17),
    (-15, 34, 13, 51, -43, -17, -8, -13, 9, 30, -32, 1, -43, -8, 3, 60, 0, -6, 16, -12, 8, 11, 4, 10, 28, 17, -13, 17, 14, 18, 20, -55, 3, 30, -22, 40, -41, -15, -65, -35, -21, 14, 1, -19, -57, 37, 26, 2, -29, 1, 30, 3, 36, 23, 24, 20, 10, 15, -34, -8, 32, 16, 50, -58, -7, -4, -22, 23, 16, -3, -68, -1, 14, 13, -8, 7, -30, 2, 26, 7, -21, 3, 24, -29, 24, 24, 31, 27, -8, -31, -14, 12, -11, 17, 23, -44, -13, -4, -13, 53, -45, -53, -42, 3, -9, -2, -7, -5, -59, 6, -1, 38, 16, -31, 56, 18, 8, 33, -17, 15, 8, -9, -47, 32, 37, 51, 3, -23, 28, 25, -13, 36, -39, -55, -16, -19, -6, 8, -9, -28, -54, 54, -23, 37, -26, -8, -4, -3, 5, 13, 10, 42, 26, -8, -35, 4, 20, 38, 39, -6, 8, 27, -15, 35, 52, -31, -29, -21, -2, -16, 28, -9, 4, 33, -3, 11, -6, 9, -52, -7, 9, 19, 19, 21, 11, 15, -11, 6, 1, 21, 20, 21, -22, -2, -1, 44, -4, -34, -37, 4, -36, -35, 3, -17, -64, -2, 25, -3, 19, -21, -5, -4, -6, 1, -1, 28, 9, -19, -64, 7, 36, 3, -6, -23, -1, -4, -32, 36, 29, -10, -4, -17, -25, -10, 34, -17, -6, 0, 7, 7, -4, -29, -42, -3, 25, -8, -1, 45, 0, -11, -62, -20, 37, 6, 20, -8, -15, 20, -26, 0, -19, -7, 20, 13, -22, -14, 37, 3, -3, 1, -13, -51, 2, -3, -18, -2, 4, -16, -12, 24, 9, 14, -22, -13, -17, 42, 32, 15, -7),
    (-17, 7, -31, -43, -11, -13, -28, 26, -25, -24, 20, -47, -21, -11, 27, -3, 15, -15, -51, -10, -19, 14, 7, 10, 24, -53, 15, 4, 12, -18, 2, -46, -47, -21, 29, -36, -51, 3, -27, 31, 3, -18, 22, 8, 30, 1, 6, -11, 44, -22, 10, -5, 22, -20, 6, 9, -26, -43, -67, -38, 2, -50, -2, 7, -30, 13, 38, -29, -29, 1, 0, 14, -6, -42, 57, -3, -20, 5, 36, -44, 33, -14, -26, -17, -25, -19, -20, -1, -49, -24, -21, -8, 13, -38, 26, 7, -35, -5, -9, 4, -27, 35, -53, 20, -50, -1, 19, 16, 20, -30, 36, -52, 40, 3, -28, -8, -24, -24, -17, -38, -12, -11, -26, 3, -34, -17, -16, 27, -16, 10, -37, 29, 32, -14, -13, 11, -40, 4, 7, -40, 2, 0, 52, -21, 48, 30, -9, 20, 0, -4, -29, 50, 0, 9, -47, -5, -33, 14, -29, -9, -31, 10, 17, 14, 2, -15, -25, 18, 11, -5, 23, -28, 0, 0, 38, 22, 2, 50, -15, 46, -26, -35, -33, 33, -13, 8, 4, -3, -26, 0, -36, 11, 25, -24, -32, -18, 23, 34, -45, -16, -34, 3, 21, -34, -6, 11, 14, 6, 11, 34, -7, 9, -36, -26, -13, -12, 15, -25, -20, -25, -45, -35, 1, 32, -10, -20, -25, 20, 7, 22, 9, 47, 26, -42, 38, -38, -27, -3, 34, -22, 56, 26, -19, -30, -2, 4, -26, -12, 22, -40, 20, -32, -14, -19, 40, 19, -38, -5, -32, 17, 30, 24, 0, -8, 16, -50, -10, -28, 32, -39, 47, 25, 20, -28, 2, -37, -34, 9, 4, 23, 0, 16, -35, -24, -29, -1, -18, -35, 7),
    (-5, -26, 3, 0, 5, 38, 41, -6, -33, 0, 5, -11, 17, 54, 14, 20, -19, -13, 28, -13, 17, -28, 25, -32, -21, 38, 47, -17, 47, 49, 23, -6, 12, -20, 10, -33, -8, 5, 28, 4, 19, 13, 27, -9, 43, 38, -11, -14, 2, 55, 14, 4, -29, -61, -32, -14, 9, -22, 38, 6, 12, 14, 34, -4, -17, 23, -42, -14, -6, -55, -22, -2, -3, -26, -15, 23, -4, 46, -43, -2, -16, 23, -14, -23, -36, -8, -10, 15, 4, -38, -20, -20, -40, -1, 14, 2, -21, -23, 11, -18, -9, -30, -24, -17, -4, -44, 39, -24, 10, 53, 24, -20, -21, -9, 0, -36, -22, -21, -21, 9, -20, -9, -17, -6, -2, 21, 21, 50, 1, -1, 31, -25, -13, 18, 17, 14, -19, 6, 10, 40, -11, 51, 5, -44, 5, -3, 21, -31, 28, -22, -25, -18, -8, 12, -6, -24, 42, 13, -30, 24, 20, 14, -19, -15, -35, 17, -7, -19, -3, -53, -31, 37, 21, 23, 0, -50, 3, -38, 25, -6, -37, 3, -4, 24, -31, -7, 13, 5, 28, -42, -28, 4, -27, 6, -19, -25, -18, 41, -11, -12, -11, 15, -28, 16, 45, 15, -25, 25, -26, -26, -15, -4, 15, -2, 29, -24, 8, -13, -14, 7, 42, -14, -32, 39, 11, 9, -31, -20, -10, 24, -38, 14, -14, -1, -32, -47, -16, -10, -11, 32, 11, -7, -31, 56, 26, -30, -9, -51, 19, 16, 15, 20, 5, -28, -3, -4, -15, 4, -11, 8, 27, 0, 7, 13, 19, -23, -22, 6, 36, -3, -33, -21, 2, -64, -26, -7, -4, 21, 3, -18, 38, 16, -21, 16, 12, 2, -30, 30, -16),
    (-19, -27, -14, 26, 14, 28, -14, -17, -27, 21, -23, -41, 13, -2, 16, 9, -23, 26, -47, 49, 25, 3, -6, -27, 36, -13, 33, -10, 14, 40, 16, 4, 25, 22, 16, 1, 41, 54, -7, -11, -24, -6, -35, -42, 20, 29, 7, -8, -45, -15, -43, 12, -14, 18, -7, -33, -3, -10, 26, 28, -7, -8, 50, 26, 13, -14, 23, -5, 5, -4, -25, -22, -23, -32, -8, -31, -21, -5, -30, 15, -10, -15, -22, -17, -20, 23, 19, -28, -2, -11, 35, 2, -15, -8, 32, -12, -23, 11, -3, 11, 46, 40, -16, -23, 26, 47, 8, 23, 32, 18, -34, -23, -1, 20, 37, 20, 26, -19, 40, -22, -1, 50, 17, -31, 0, 12, 41, -1, -37, -5, 13, -25, 43, 9, 7, -3, 1, 40, -28, 11, 2, 48, 5, -27, -17, 44, 11, 13, 23, -2, 44, -46, -27, 6, 1, -10, 13, 24, 41, -32, -22, -15, -3, -23, 15, 15, -20, 24, 12, 17, -13, -34, -1, -6, -24, 34, -20, -1, 46, 0, -25, -18, -7, -10, -9, -3, 19, 28, -27, 19, -2, -24, -39, -6, -16, -51, 9, -33, -28, -42, -32, -1, -32, 2, -25, 34, 13, -47, 23, -11, 21, 26, 23, 10, 12, 23, 6, -20, -19, 17, 14, -27, 16, -9, -28, 31, -10, -34, -26, 10, 31, 12, -16, -4, 18, -3, -4, 7, -1, -30, -3, -8, 22, 30, -17, 9, 11, -47, -32, 16, 20, -5, 18, 18, -4, -5, 7, -9, -30, 13, -19, 19, -9, 7, 27, 37, 0, 33, 9, 38, 14, -36, 2, 19, 48, 31, 3, -40, 48, -44, -5, -15, -17, -19, 46, 17, 32, -9, -5),
    (13, 25, 6, -8, -27, -26, -45, 2, -13, 34, 7, 25, 17, -4, 7, 19, -23, -16, -43, 34, -5, 20, 18, -4, -12, -24, 19, 4, -4, -25, 33, 15, -1, -13, -9, -38, -16, -6, 0, 34, 21, -19, 15, 22, 34, -12, 5, -11, 17, 14, -56, 26, 17, -14, 20, -33, 13, -3, 34, -18, -17, 2, 17, 12, 18, -49, 16, -22, -5, 17, 32, 13, -8, -7, 27, 12, 29, -7, 1, 9, -23, 3, -19, 1, 16, 8, 27, 24, -21, 3, 24, -9, 19, 9, 16, 44, -40, -45, 22, 2, -21, 43, -33, -29, -12, -1, 16, -6, -15, -15, 9, 21, -4, 6, -70, 47, -30, -41, 31, -23, -24, -3, 27, -30, 16, 17, 0, 7, -22, -30, -6, -35, 34, -12, 28, 44, -39, -7, 7, -20, 54, -3, -7, 13, -7, 12, -61, 28, -5, 3, 12, -31, -26, -16, 34, -8, -8, -34, 30, 50, 4, -21, 11, -15, 5, -6, 23, 28, -2, -33, -16, 8, 9, 6, 7, -10, 19, -2, 12, -13, -1, 1, -18, 8, -15, -17, -4, -24, -28, 24, 17, 3, -10, -39, 8, -16, 45, 20, -16, 34, 20, -12, -11, 25, 23, -28, 9, -15, -31, 14, -22, 61, 28, -18, 11, -19, -22, 25, 38, 14, 17, 17, 39, 23, 18, -16, -18, -26, 58, 11, -8, 5, -28, 31, 9, 20, 19, -19, 2, -11, 13, 21, -28, 60, -33, -14, -12, -1, 0, 31, 27, 17, -42, -9, 15, -11, 7, -33, 23, -21, 8, -9, 31, 38, -10, -2, 21, 13, 9, -5, -1, -18, 4, 20, 42, 7, 5, -9, -19, 27, -6, 14, 7, 37, -17, 16, -19, 22, 13),
    (-18, 24, 1, 11, -44, 16, 8, 11, -21, -50, -12, 14, 6, 20, 21, -17, 6, -4, -4, -34, 14, 0, 20, 18, -23, -23, -25, -24, -15, -40, 29, -13, -6, 27, -33, -17, -20, 5, -52, 16, -43, -37, -3, -7, -1, 5, 27, -35, 8, 3, 2, -30, -26, 11, -1, 18, -24, -75, 0, -5, -26, -36, -2, 27, -19, 11, -18, -33, -16, 12, -34, 22, -30, -41, 25, -20, -3, 19, 29, -8, 12, -4, -3, -19, 23, 41, 19, -24, -27, -56, 11, -39, 2, -21, -11, 8, -10, 43, -2, 3, 15, -20, -27, 6, -53, 27, 0, 25, -2, 15, 2, 24, -3, -30, 46, -31, 26, 22, 8, 28, 7, 3, 42, -16, -14, 32, -5, 17, -7, 29, -24, -4, 37, 14, -42, -23, -8, 2, 12, 6, -18, 21, -17, -28, -13, -3, 17, -52, 21, 43, 38, 15, -18, -33, -5, -46, -12, 56, 23, 17, 20, 32, -5, 32, 39, 17, -21, -6, -28, -17, -36, 19, -14, -15, -30, 6, -16, -28, -16, -1, 14, 55, 29, 32, -8, -43, -9, -32, 8, 32, 59, 5, 10, -23, -14, 33, 19, -1, 5, -24, -2, 28, 16, 47, 19, 24, -54, 26, 4, -3, 47, 1, -10, 5, 9, -10, -21, 9, 38, 1, -20, 68, 32, 22, 17, -10, -13, 14, 1, 15, -31, 6, -50, 31, 4, 61, -26, -3, -52, 5, 20, -2, 28, -51, -16, 34, 5, 24, 19, 17, 19, -45, 9, 48, 19, 0, -21, -26, 0, 36, 4, -29, 12, 8, -45, 24, -40, 36, 21, 3, -10, -49, 6, -16, -18, -29, 22, 51, -2, 8, 18, 2, -5, -33, -11, 15, 18, 2, 1),
    (9, -7, -28, -32, -44, 11, -30, 31, -7, -20, -10, 0, -6, 7, -30, 3, 26, 1, -49, -1, 7, -7, -34, -31, -19, -22, 10, 10, 3, -39, -54, -32, -18, -32, -48, 9, -2, -21, -39, 58, -28, -44, -12, 15, -7, -36, -17, 17, 20, 3, -18, 40, -54, -25, -34, 13, -12, -3, 6, -14, -17, 6, -46, -8, -55, -12, -1, 33, -1, -11, 33, 27, -16, -55, 11, 13, -13, -7, -10, -32, 13, 23, -24, 15, -12, -2, -40, -4, -6, 3, -10, -15, -28, -33, -18, 24, -45, -13, -7, -8, 24, -19, 12, 14, -18, -26, 44, 1, -20, -40, 17, 14, -20, 13, 30, 11, -40, -8, -23, -1, -25, 10, -27, 1, -16, 18, 20, -40, -21, 11, -25, -20, 49, 25, -6, 18, 40, -7, 4, -6, -42, -44, -17, 4, 4, 9, 2, 9, -17, -30, 3, 6, 35, -4, 36, 1, -16, -32, -7, -17, 4, -1, 16, -20, 13, -16, -1, 40, 22, -11, 6, -16, -16, -16, 21, 24, 33, 17, -24, 14, -21, -3, 24, -2, 14, 19, -19, 16, -33, 18, 20, -1, 1, -7, -11, 23, 34, 11, -27, 21, 26, 9, 33, 16, 7, -41, -6, 45, 18, 1, 48, 3, -5, -14, -42, 8, 42, 13, -17, 9, 12, -20, -33, -43, 8, -2, 36, -16, 27, -6, 6, 24, 12, 3, 12, -21, -1, -11, 16, 56, -16, -22, 43, -21, 17, -17, -7, 50, 12, 23, -14, 8, 18, -11, -13, -37, 23, 1, -6, -12, 26, -27, -26, -25, 39, 32, -33, -24, -11, 7, -26, 23, -16, -5, 7, 25, 27, -44, 13, 13, 1, -17, 52, -7, -31, 12, -12, -1, -12),
    (-7, -20, -2, -7, -10, 1, 32, -11, 24, -2, -2, -12, 2, -24, 5, -7, 18, 18, -10, -19, 9, 13, -10, -7, -14, -33, -32, -14, -23, 7, 34, -22, -23, 40, 39, 20, -39, -29, 20, -23, 26, 25, -60, -23, -29, -27, 3, 14, 27, 2, 37, -39, 14, -38, -17, 18, 28, -62, 53, -28, -18, 22, -7, -61, -16, 18, 0, 18, -32, -39, -13, -64, 20, 27, -50, -24, -43, 17, -5, 0, 6, -13, -4, -41, -33, -20, -27, 21, 28, -43, 14, -43, -10, -23, -13, -32, -9, 21, 18, -10, -4, 29, -13, -20, 45, -10, -64, 1, 18, -29, -50, 37, -2, 7, 30, -2, -4, 20, -29, 23, 7, -20, 5, -2, 13, 24, -11, -8, -9, 19, 5, -30, -54, 38, 23, -47, 25, 10, -101, -17, -8, -3, 10, -34, 18, 3, 40, 1, -44, 15, 3, -40, -1, -56, -1, 4, 35, 0, 4, -64, -33, 12, 33, 13, -26, -22, -15, -12, 27, 24, -79, -26, -39, -15, 28, 1, -2, -69, -3, -41, -36, 24, -5, -18, 42, -47, 13, 31, 46, 4, 0, -17, 10, -4, 23, 19, -45, -38, 14, 25, 10, -19, -43, 29, -25, -25, -23, 20, -26, 16, -7, 3, -37, 26, 9, -8, 9, -9, 15, 25, -6, -9, 20, 8, 0, -21, -42, -10, -49, -11, 12, -3, -12, 50, -41, 23, -8, -13, 23, -16, -3, -13, -8, -7, 15, 27, 23, 3, -1, -19, -33, 20, 48, 21, -4, -30, -30, -37, 1, 0, -17, 7, -44, -28, -30, 24, 9, 3, -19, -20, 33, 17, 9, -72, 31, -14, -24, 6, 21, -27, 34, -25, -13, 8, -11, 5, -14, 12, -6),
    (1, 21, 10, 52, 0, -32, -4, -44, 10, 4, -7, 28, 13, 3, -17, 47, -10, -21, 57, 10, -40, 34, 2, -8, -21, 20, 25, -2, -8, 39, -28, -10, 18, -5, -47, 20, -30, 16, 43, -14, 26, 11, 3, -6, -16, 16, -38, 14, 16, -1, 52, -16, -27, 12, 42, -33, -40, -20, 41, -32, -18, 0, 18, -4, -12, 32, 13, 13, -2, -3, 32, 26, -13, -14, 20, -11, 32, -15, 21, 5, -4, -30, 3, 28, -39, 10, -11, -21, -32, -12, 20, 7, 17, 24, -8, -41, -12, 0, 49, -17, -22, -6, -16, -10, 11, -24, 5, -8, -3, -27, -50, 7, 15, -53, 27, -37, 23, -19, 7, -10, -19, 8, -25, -50, 2, -47, -46, -21, -4, -38, -6, -2, -5, 34, -36, -6, -35, 1, -9, 40, -39, 2, -6, 6, 20, -60, -40, 21, 25, 22, 37, -4, -11, -13, 24, -34, 16, -21, -44, -48, -26, 9, 1, -9, 4, 22, -60, -3, 11, -31, 12, -21, -45, 2, 0, -1, -62, -20, -28, 10, -11, -13, 3, -32, -5, 0, 16, -33, 2, 22, -45, 7, 37, -10, 21, 30, -33, 28, -43, -24, -2, -36, -10, 16, 7, -55, 1, -8, 49, -35, -18, 27, 7, 14, 40, 11, 33, 6, -34, -24, 11, -34, -12, -25, -8, -28, -13, -5, 6, 18, -30, -28, -29, -37, -34, 4, -14, -1, -2, 29, -4, -23, -38, -9, -6, -43, 40, -33, 34, -38, 18, 12, 19, 32, -33, -7, 2, -47, -10, 7, 4, 9, -32, 45, -42, -5, -20, -22, -8, 16, 9, -1, -35, -26, -27, 26, -7, 9, -8, -23, 12, -21, -44, -2, 19, 13, -13, 11, 6),
    (-5, -21, -7, -42, -26, -56, -3, 42, -20, 0, -1, 22, 18, 39, 38, -22, 25, -24, 9, -21, 7, -2, 10, -5, 18, 30, 11, -3, -35, 32, -4, 23, -13, 4, 1, -11, -40, -6, 1, 30, 15, 6, 48, -47, -10, -20, 33, -6, 10, 9, 6, -4, 38, -25, 45, 2, -16, 41, 27, 8, 15, 33, 32, -23, 15, -34, -9, -15, -26, -11, 4, -27, -13, -11, 29, 17, 14, 11, 30, -45, 33, 5, -26, -14, -8, -33, 42, 0, 6, 38, -13, 50, -22, -21, 12, -36, -47, -25, -23, -40, -31, 3, -5, -14, 32, -95, 41, -26, -48, 4, 65, -28, 41, 8, 6, -9, 11, -14, -48, -6, -22, -30, 2, 27, 5, -39, 12, 27, -60, 12, -33, 39, -25, 21, -37, 11, 1, -36, 44, -9, -46, 21, 47, 33, -2, 10, -39, -24, -7, -30, -4, -9, -28, -45, -26, 35, 8, -37, -9, 11, -35, -35, -31, 12, -8, 22, -20, 1, 25, -39, 29, -28, -12, -22, 62, 1, 4, 55, -3, 17, 5, -14, -34, -22, -1, -18, 5, 25, -13, -43, 14, 40, 25, 29, -7, 12, 42, 27, -11, -1, 25, 9, 31, 17, -5, 21, 29, 9, -28, -1, 23, -39, -24, -35, -35, 9, -6, 24, -7, 4, 10, -5, 8, -8, -18, 38, -28, -29, 9, -13, 14, -17, -15, 5, 6, 13, -27, -38, 13, -12, 13, 25, -3, -25, 7, -10, 4, -22, 4, 21, -32, -37, -23, -6, -27, -1, -29, -6, -4, -40, -6, -9, 38, 26, 21, -14, 17, -8, 8, 14, 10, -8, -36, 21, 8, -43, 37, 38, 21, 36, -2, -13, 14, -38, -34, -1, 12, -3, 36),
    (-10, 20, -8, -36, -15, 36, 11, -33, -7, 13, -33, -2, 8, -17, -18, 37, -28, -48, -39, -18, -34, 17, 28, -38, 0, 24, 38, 2, -5, 34, 30, 8, -20, -15, 6, 4, -14, 58, 15, -35, -20, 30, -3, -14, 19, -1, 30, -2, 21, -35, 42, -36, -10, 49, -16, -21, 10, 44, -37, -25, 30, -23, -16, 42, 16, 18, 1, -38, -47, 37, -16, -19, -6, 4, 8, 14, -50, -19, -7, -28, -8, 1, 46, -32, 3, 72, -37, -16, -15, 18, -76, -13, -30, 2, 19, 5, 4, 37, 0, 4, -35, 0, 12, 29, 8, 34, -29, 10, -18, 21, 58, -9, -32, -19, -20, -11, -10, 57, -6, -23, -22, 38, -26, 45, 9, -3, -19, 16, 39, 34, 4, -27, -34, 25, 0, -33, -17, -9, -41, -22, -47, 19, 37, -2, -30, -47, 48, -29, -27, 95, -2, -24, 6, 8, -45, 29, -7, -20, -37, 37, 34, -11, 30, 21, -25, 46, -27, -22, -25, -6, -8, -42, -40, -27, 4, 26, -5, -38, 20, 23, -21, 41, 12, 21, 16, 22, -3, 4, 25, -48, -45, 26, 23, -10, 24, -14, -41, -20, -19, 1, 12, 16, -5, -10, 14, -24, 42, -17, 18, -7, 3, 14, 31, 42, 2, 30, -7, 31, -35, -11, 37, -56, -20, -10, -9, 16, 38, 13, -21, -1, 10, 14, 39, 37, -45, 19, -33, -29, 24, 27, -21, -9, -21, -6, 20, 21, -26, 14, 9, 31, -30, 15, -7, -28, -29, 2, 0, -14, 23, -18, -1, -12, -21, -26, 19, -7, -4, -23, -3, 0, 8, 21, -5, -14, -22, 23, -38, 23, 30, -21, 16, 2, -5, -25, 21, -33, -29, 27, 2)
  );
  ----------------
  CONSTANT Layer_8_Columns    : NATURAL := 4;
  CONSTANT Layer_8_Rows       : NATURAL := 4;
  CONSTANT Layer_8_Strides    : NATURAL := 1;
  CONSTANT Layer_8_Activation : Activation_T := relu;
  CONSTANT Layer_8_Padding    : Padding_T := same;
  CONSTANT Layer_8_Values     : NATURAL := 48;
  CONSTANT Layer_8_Filter_X   : NATURAL := 3;
  CONSTANT Layer_8_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_8_Filters    : NATURAL := 48;
  CONSTANT Layer_8_Inputs     : NATURAL := 433;
  CONSTANT Layer_8_Out_Offset : INTEGER := 3;
  CONSTANT Layer_8_Offset     : INTEGER := -1;
  CONSTANT Layer_8 : CNN_Weights_T(0 to Layer_8_Filters-1, 0 to Layer_8_Inputs-1) :=
  (
    (18, -31, -9, -9, 15, -24, 34, -19, 24, 27, 6, -9, 17, -24, -18, 17, -2, -7, -8, -30, -7, -10, -26, -20, 31, -15, -5, -7, 9, -27, 11, 11, -26, 11, -7, -1, 35, -9, 13, 11, -1, 23, -27, -30, 9, 11, -10, -42, -3, -36, -25, 14, 12, -3, 16, -7, -8, 25, -7, 17, -5, -17, -21, 28, 14, 6, -14, -12, -7, -16, -24, -17, 26, 0, -12, 46, 19, 3, -19, 7, 2, 15, -19, -10, 21, -26, 63, -26, 1, 3, -51, 8, -17, 1, 18, -4, -18, 17, -37, 17, 7, 17, 15, -10, 45, 33, -16, -6, -6, -38, -22, 35, -25, 26, 23, -13, 14, -33, -13, -18, 38, -4, 17, 36, 24, -1, 3, 13, -1, 0, -22, 1, 26, -5, 16, 10, 3, 33, -27, -10, -1, 22, -15, 25, 9, -10, -26, -24, 0, -35, 38, -20, -2, 4, -13, 32, -4, -22, -14, 30, -22, -10, -30, 0, 41, 26, -31, -6, 22, 7, -17, 7, 17, 0, 2, 11, 13, -14, -9, -15, 26, 3, -28, -30, -7, -14, 2, -9, 9, 11, -26, -10, 17, 16, -1, -4, 23, -4, 18, 15, -15, -11, -7, 4, -10, -6, -32, 7, 44, 19, -18, 25, 25, -14, -65, 3, 1, 31, 26, 27, 10, -25, -14, -26, -15, -25, 17, -28, 13, -13, -16, -5, 9, 9, 0, -26, 37, -3, -38, -21, 22, 14, 16, -18, -15, 19, 35, -39, -1, -10, 3, -20, 18, -7, -22, 27, -12, 17, 1, 21, -1, -32, -41, 27, -14, 16, 35, 22, -14, 7, 21, 12, 21, -29, -13, 17, 23, 1, -17, 15, 17, 34, 20, 20, -14, 28, -38, -17, 6, -25, 30, -41, 0, 17, 19, -44, -16, 14, -50, 17, -14, -35, -23, 5, -5, 1, 0, 12, 18, 22, -22, -22, -4, 5, 19, 29, -35, -31, -23, -3, 8, -22, 9, -23, 8, 14, -9, 8, 18, -9, 42, -24, 9, -20, -3, 3, 5, -21, -54, -60, -14, 42, 34, -31, -6, -16, 39, 6, 11, -3, 1, 13, -45, 15, -27, 1, -12, 25, -32, -20, -22, -4, 30, -13, -17, 4, -15, -11, -6, -43, 6, -13, 10, -22, 12, 27, 1, 17, -16, 5, 20, -5, -1, 34, 22, -37, -13, -29, -18, 56, -12, -72, -17, 30, 1, -7, 30, -4, 22, -9, -25, -23, 33, -4, 42, 21, -42, 14, 11, 20, 6, 10, 5, -20, -15, 27, 4, -41, 4, 9, 26, -48, -35, 8, 38, 13, -39, 4, 7, 11, -37, -13, -6),
    (-14, -12, -27, -47, 15, -9, 20, 8, 30, 16, -1, -9, -11, -8, 6, 32, -31, -34, -27, 23, 18, -1, 35, -31, -33, -20, 25, -6, 21, -20, -38, -15, 14, 7, 7, 32, 34, -29, -7, -7, 22, 9, 37, 14, -17, -38, 15, 13, -17, 1, 3, -21, 19, 7, -12, 0, 26, 3, -21, -34, -18, -8, -13, -13, -4, 16, -29, 26, -14, 32, -14, 22, -12, -15, 15, 11, 36, -10, -22, 6, 20, 19, 29, 12, 6, 0, -17, -3, -30, -12, 28, 10, -25, -6, -12, -5, -35, -3, -7, -4, 0, 18, 2, 6, 7, 4, -42, 1, -25, 18, 34, 10, 4, -2, 12, 11, -12, 20, 0, -15, 22, -42, 3, -35, 10, -13, -12, -12, -16, 47, 3, -10, -16, 25, -32, 36, -15, -27, 16, 10, -48, -22, 18, 24, -31, 21, 14, -12, -16, 18, -11, 9, -6, 2, -15, -18, -23, -48, -39, -6, 16, 12, -16, -39, -19, -19, 66, 18, 13, -13, 20, -3, -2, 11, 30, -29, 3, 12, 26, 20, -40, 51, -15, 4, -8, -23, 58, -23, -6, -50, 26, 3, -33, -5, 2, 5, 6, 17, 1, 35, -6, 2, -35, -16, -2, -29, 12, -23, 44, 31, -21, 3, -50, 7, 20, 18, 45, -12, 20, 43, 30, -29, -41, -29, -49, -18, -5, -17, -5, 34, -8, -30, -9, -2, 27, -15, -12, -17, 10, 17, -14, 20, 38, 16, -22, 21, 26, 48, 25, 39, -34, 3, 4, -16, 9, 32, 15, -4, 1, 11, -31, -46, -16, -30, 13, -13, 27, 30, -8, -11, -8, 19, -5, -8, -24, -25, -13, -9, -29, 16, -16, -5, 28, -41, -41, 25, 16, 17, 23, -16, 31, -16, -11, 25, 19, -13, 8, -12, 11, -3, -6, 3, -25, 5, 22, 14, -13, 3, -7, -15, 13, -17, 2, -7, -11, 35, -1, -12, -10, -3, -8, 2, 6, 26, 7, 28, 12, -14, -15, 8, 7, -51, -36, -5, -13, -16, -25, 14, -8, -16, -2, 8, 11, 23, -12, 14, -1, -2, -1, 6, -9, 7, 4, 6, -12, 16, 5, -8, 19, -23, -14, -12, 33, 25, -16, -16, 26, -4, -24, -7, 7, -34, 21, -13, -14, 5, 18, 9, -16, 26, -18, -18, 10, 8, 16, -28, -17, -23, -22, -28, -5, -7, -36, 8, 8, -48, -5, 40, -14, -17, -62, 17, -9, -2, 32, 23, 2, 6, 3, -25, -8, -18, 3, 17, -18, -15, -10, -26, 8, -17, -14, 0, 4, -41, 15, -13, 33, 2, 9, 20, 8, 30, -5),
    (-27, 32, 9, 51, 15, 42, 8, -9, 2, -6, -14, -4, -32, -28, 9, 33, 24, 34, -26, 6, -28, -12, -7, 1, -10, -23, -15, -17, -3, -19, 21, -6, -9, -18, -6, 10, 12, -9, 7, 38, 41, 28, 14, 12, -13, -8, 0, -28, 5, 22, 6, 28, 30, 19, 4, -21, 27, 9, -2, -14, -7, -44, -7, 30, -1, 20, 8, -25, 0, 38, 17, -3, 5, -9, 43, -17, 14, -39, -23, 21, -10, 15, -11, -6, 19, -17, 5, 7, 18, 20, -13, 26, 18, -8, 15, 13, 0, 25, 19, -11, -4, -26, -20, 4, 22, -11, 9, 13, -48, -21, 5, 6, -12, -51, 13, -12, -7, 22, 5, 21, 1, 4, -3, -16, 8, -20, 10, -6, -1, 26, -20, 3, 18, -29, -36, 18, 34, 23, 31, 20, -35, -35, 15, -27, 11, 20, 12, -1, -9, 35, -5, -28, 30, 11, 8, -17, -38, -12, -28, -7, -31, 23, 1, -8, -29, -32, 22, 28, 15, -7, -17, 1, -40, 9, 2, 29, 2, -7, -28, -11, -10, -5, -14, -26, -19, 14, -39, 36, -1, -11, -20, -10, 11, 15, 25, 16, -12, 2, -11, -14, 0, 0, 40, -33, 16, -38, 30, -11, 0, -15, 22, 25, -27, -18, 8, 3, 25, -30, -2, -14, -55, -14, 35, 24, 10, -1, -5, -7, 31, 1, 13, -26, -22, -36, -38, 25, -32, 0, 43, 42, -27, 28, 4, 4, -16, -38, -9, 24, -3, -19, 11, -7, -7, -7, 3, 37, 21, -17, -18, 15, -39, -26, 21, -24, 8, -21, 32, 4, -41, -13, -14, -4, -12, -20, -3, -5, -10, -20, -3, -21, -23, -7, 11, -5, 16, 10, 10, -11, -13, -11, 17, 23, -4, 2, -2, 25, 35, -36, -45, -31, -44, -25, 16, 42, 5, -19, -16, 9, 7, 21, -12, 2, -27, -3, -3, 0, 16, -9, 11, -48, 17, 14, -14, 22, -35, 10, 18, -30, 11, 14, 22, 4, 9, 13, 2, -9, -29, -20, -17, -7, -2, -29, -6, 9, -22, 0, -9, 10, 4, 20, 20, 4, 4, -8, 3, -31, 11, 28, 3, -22, -35, -39, 0, 1, 30, 24, 55, -29, -25, -30, -8, 14, -38, 32, 7, -32, -33, -24, 8, 29, 12, -20, -7, 22, -6, 18, 8, -23, -12, -27, 6, -26, -29, -1, -1, 6, 6, 19, 0, -20, -2, 5, 16, -23, 22, -1, -25, -24, -21, -16, -18, -26, -7, 30, -15, 4, 18, 2, 23, -17, -5, 3, -5, -22, 15, 3, -27, -9, -17, 24, -13, -24, 7),
    (-8, -27, 0, 15, 24, -10, 13, 42, -13, -49, -42, 66, 8, 5, 28, -38, 40, -9, 2, -8, 25, 29, -25, 17, -2, -22, -49, 19, -5, -14, 5, 3, 7, 18, 12, 28, -16, -5, 12, -16, -7, -42, -48, 24, -37, -9, 15, 1, 3, 14, 17, -21, -11, 10, -8, 35, 14, 7, 3, 7, -9, 4, 6, -2, 7, 0, 21, -15, -15, 16, -38, -9, 39, -25, -10, -24, -7, -9, -26, 4, -31, -6, 13, -3, -15, -8, 25, 14, 14, -1, 6, 7, -17, -5, 15, -10, -8, 3, 21, -41, 7, -6, 36, 5, 16, 24, -20, 20, 43, 1, 18, -7, -3, -30, 10, -31, -37, 23, -8, -2, 23, 25, 5, -17, -9, -19, -24, 0, 24, -11, -11, 22, -6, 17, -36, 32, 17, -17, -14, -7, 6, 26, -36, 8, -22, 13, 64, -33, -7, -3, 0, 9, 10, 1, 1, -11, 2, -16, -23, -7, 16, 6, -9, -21, -38, -22, -30, 16, 26, 2, 18, 3, -2, 35, -6, 11, 7, -8, 5, 21, -39, 24, 31, 18, -25, -13, 22, -28, -4, -18, -14, -49, -26, 1, 55, -40, 15, 1, 35, 23, 16, -6, -25, -12, 44, 0, 17, -3, -31, 2, 7, -7, 14, -14, -5, 11, 11, -8, 3, -14, -10, 3, -22, -7, 10, -31, 18, -21, -1, 47, -17, 30, -1, -1, 37, 3, -15, 21, -46, -16, 24, -32, -17, -31, -41, 2, 35, -41, -11, -10, 10, -18, -11, -9, -22, 26, -20, 2, -22, 25, 18, 14, -51, -5, 2, -4, 30, 12, 13, -5, -16, -33, 27, -3, -1, 25, -7, 0, 1, 28, 11, 13, 1, 10, 2, 30, 1, 24, -1, 11, -3, 0, 18, -2, 10, 34, 10, -1, 9, 6, 5, 30, 19, 20, -42, 9, -19, -2, -16, -4, 17, -21, 14, 23, 47, 19, -7, -20, -44, -15, 12, -33, 7, 12, 17, -4, -9, 31, -9, 6, 0, -6, -20, -23, 13, -30, -9, -18, 22, -26, 7, 38, -21, 16, -32, 26, -13, -43, 10, 16, -14, 21, 14, 24, -7, -22, -23, -12, 25, 31, -16, 28, 22, -16, -11, -7, -28, 22, 19, -2, 18, 31, 13, -5, -37, -29, 22, 3, 32, 15, 23, 40, -14, -21, -3, -20, 4, -13, -23, -2, -16, -7, 8, -8, 1, 5, 17, -29, -32, 19, -14, 12, -29, 17, -2, 25, -34, -2, -9, -10, -5, -16, -6, -23, -15, -8, 14, -13, 3, 43, -14, -21, -12, -12, 8, 35, 28, -23, 16, -1, -21, 14, -2),
    (-30, 18, 16, 15, 19, 20, -40, -8, -6, 21, -16, 6, -12, 33, -26, -15, 7, -12, -4, 22, -44, -19, -26, 0, -3, -26, -3, 14, -9, -12, 2, 28, 13, -8, 15, 22, -12, 6, 12, 4, -20, 2, -6, 30, -3, 7, 15, 23, -13, 28, -18, -1, -15, 22, 17, -18, -5, 11, -20, 7, 24, 4, 24, 2, 13, 36, -21, -3, -14, -29, -47, 30, -35, 4, 2, -6, -2, -33, -3, 13, 6, -3, 16, 2, 21, -30, 13, 19, -19, 45, -24, -3, -38, 1, -9, 16, 3, -12, -15, -56, -10, -2, 20, -12, -2, -32, -6, 19, 17, 28, 12, 32, -8, 18, 0, 32, -3, -15, -17, 11, -12, 8, -44, 27, 16, -42, -35, -4, -4, -4, -2, -10, 25, 15, 1, 4, -16, -2, -13, 12, -2, 21, 11, 33, -8, 19, 4, 31, -8, 8, -53, 5, -1, -22, 10, -1, 25, 23, -27, -14, 11, -5, 14, 22, -33, 9, 15, 20, -26, -17, -35, -14, -15, -19, -15, -23, 9, 0, -3, 0, -27, -23, 15, -19, -43, -13, -17, 12, -48, 18, 8, 34, -29, 18, -9, -7, 4, 15, -32, 12, -10, 5, -13, -22, -27, 28, 3, 8, 6, -3, -14, -37, -6, 15, -5, 35, -21, -44, 7, -6, -14, 1, 2, -25, -29, -1, 3, 8, -5, -18, -53, -35, 6, 35, -5, -1, -33, -1, 8, 27, 9, 4, -31, 21, 14, -8, 10, 25, 20, -22, 13, 1, -3, 26, 38, 8, 1, 1, -12, 21, 39, 7, -16, 21, -9, -17, -19, -9, 3, -34, -21, -8, 7, 9, -34, -24, 14, 23, 0, -4, -7, 7, -19, 18, 6, -3, -6, 6, -39, 58, 21, 67, -20, -37, -30, 52, 8, 29, -48, -21, 1, 0, -33, -12, 26, 10, -3, -36, -81, -36, 9, 2, 28, -5, -31, 22, -4, -5, 0, -28, 5, -2, 3, 0, -40, -30, 32, -24, -6, 3, -52, -48, 0, -7, 40, 5, 18, 48, -6, 42, -18, 2, -20, 24, 8, 38, 3, -51, 3, -10, 16, 20, -17, 0, 11, -13, -47, -46, -31, 3, 13, -11, -9, 40, -4, -8, -28, -22, -1, 14, -1, 4, 5, -7, -19, 2, 3, -32, -6, -25, 12, -5, 35, -14, -8, 16, 32, 22, 4, -13, 7, 49, -2, 15, -18, -45, 35, -23, 3, -19, -13, 15, 8, 9, -5, -22, -7, 11, 17, -8, 17, 35, 9, -23, 55, 5, 12, 20, -25, -7, -6, -13, 33, 0, 9, 6, 17, 11, 4, -20, 40, 18, 12),
    (-5, 23, -44, -43, -22, 12, -52, -6, 10, -20, 6, -14, -22, 29, 7, -17, -15, -34, 37, -2, -26, -1, 19, 35, -18, 3, -48, -28, 14, 4, 9, 3, -31, -5, 8, 27, -6, -3, -14, -55, -12, -33, -30, -8, 1, 7, 13, 36, -16, 41, -17, -34, 30, 27, -17, 6, 11, -11, -25, -3, 20, 35, 27, -28, 0, 8, 13, -23, -6, 15, -3, -5, 4, 24, -79, -34, 13, -29, 6, 9, 13, 12, -18, 4, 13, 20, 12, -24, -48, -4, -4, 28, -26, 18, 7, 26, -34, 43, -11, -5, -8, 26, -35, -37, -26, -1, -25, -41, 7, -8, 28, -4, 37, 43, -29, 40, -7, -12, 3, 32, -47, 2, -17, -28, 9, -21, 10, -12, 15, 39, -37, 24, 13, 28, -27, -26, -25, -24, -2, -10, -23, 5, 1, 14, 16, 10, 23, -48, 34, -33, 12, -23, 8, -1, -31, 27, 27, 36, -27, -29, 30, -46, -9, 12, -34, -13, 13, -10, -21, 2, -42, 4, -9, -8, 20, 26, 6, -11, 13, 14, -45, -14, 36, 30, -2, 0, -12, 0, 1, 17, 10, -35, -23, 15, -5, -23, 21, -20, -20, 24, 12, -15, -45, -26, 8, 15, -6, -32, 4, -52, -8, -16, 20, -12, 13, -5, 16, 26, -44, -16, -13, -12, 7, 16, 16, -17, -3, -34, -7, 32, 9, 18, 10, -11, -29, -13, -24, -6, -19, -38, -46, 44, -14, 0, -1, -7, -42, 23, -24, -13, 20, 19, 8, 8, -18, -46, 18, -37, -3, -12, 11, -11, 15, 16, 4, 6, -58, -20, 21, -17, 31, -13, -4, 27, 18, 19, -14, -29, -9, -28, -40, 43, -23, -20, -13, -1, 3, 4, 4, 17, 33, -9, -27, 36, -9, -5, -20, 4, -22, -11, -31, -9, 23, 0, 19, -33, 1, 6, 6, -18, -19, -5, -34, 6, -4, 24, -16, -4, -17, 0, 4, -13, -29, 31, -12, -29, 15, 18, -11, -20, 28, 4, -4, 21, 45, 3, -11, 29, 17, -22, 13, 10, -14, 2, -29, -24, -22, -7, 20, 18, 0, 39, -10, 11, -15, 4, -26, -17, -2, 9, -37, -1, 30, 10, 5, -6, 14, -13, 4, 8, -8, 45, 3, -6, 11, 3, 24, 23, 20, -18, 20, 17, 19, -46, 7, 20, -18, -15, -25, -43, 8, 8, -14, -25, -28, -16, 28, 11, -20, 10, 19, 3, -19, 22, -10, 38, -1, -25, -41, 28, -18, 4, 14, -13, 1, -17, -13, -40, -3, 64, -15, -28, -30, 7, 9, 15, 2, 4, -13, 7, -4, -35, 23),
    (29, -35, -14, -43, -5, -5, 10, 18, -22, -29, 10, 17, -4, -32, -7, -7, 17, 23, 26, -5, 0, -38, -18, 6, 11, 17, -6, -23, 7, -13, 6, -1, -1, -2, 12, 1, -14, 45, 7, -4, -24, -17, -15, 1, 16, -12, 13, 20, 11, 31, 12, -17, 34, 29, 29, 26, 13, 12, -7, 29, -15, -25, -15, 12, 21, -7, -3, -16, -12, -14, -3, -26, 22, 8, 34, 27, 0, -4, 13, -15, 15, 16, -11, -20, -11, 13, 18, 7, 18, 14, 7, 4, 26, -18, 14, 10, -41, -32, -2, -12, -17, -25, -10, -55, -16, -4, -16, 8, -29, -10, -14, -32, 22, -34, 18, 6, -23, -7, 41, -26, 13, -21, -14, -30, -4, -2, -10, 21, -1, 5, 12, 15, 17, 50, -20, 13, -5, 4, -26, -28, 7, -5, 18, -2, -9, 10, 18, -34, -5, -19, 5, -24, 4, -36, -13, 20, -27, -11, 23, 4, 9, -8, -4, 5, 35, 10, 26, 15, -14, 29, -20, 15, -9, -8, -43, -28, -12, 0, -16, -36, 2, -6, -36, 8, -33, -14, -26, 6, 23, 9, -32, 13, -2, 11, -23, -9, 7, 39, 18, -35, -5, -2, -19, 4, 7, -1, 25, 7, 7, -5, -59, 8, -9, 1, 45, -32, -39, 36, -24, 12, -17, 22, 7, -15, 27, 23, 10, 23, 23, 4, -7, -11, 24, -34, 36, 0, -20, 11, 7, 18, 4, 7, 4, -16, -31, 30, -24, -22, -4, -39, 20, -20, -10, 17, -2, 13, 20, 37, -23, 10, 14, 11, 7, 18, -37, -16, 24, -5, -6, -8, 19, -18, -25, -3, -36, -10, 27, -25, 17, -2, -20, -20, -11, 16, 17, -28, -5, -3, -15, 42, 17, 29, 21, 34, 7, 38, -11, 5, -23, 2, 23, 0, 30, -1, 21, -26, -45, -3, -39, -33, -8, -10, 53, -4, -7, -7, -44, -7, -25, 28, -8, 25, -29, -22, 30, -16, 0, -29, 4, -41, -19, -29, -4, -19, 16, -29, -29, 32, 42, -50, 24, -35, 18, 29, 37, -1, 1, -11, 27, -38, 2, 9, -13, 12, -40, -16, -17, -3, 15, 29, 17, -1, -1, 3, -12, -13, 13, -17, -9, 14, 6, -16, 33, 29, -28, -3, -35, -12, 10, -38, 19, -40, -7, -16, -9, 28, 17, 6, 27, 6, 34, 23, -2, 34, 23, -2, -12, -28, 20, -13, 13, -25, 18, 37, 14, -1, -22, 18, 28, -7, 8, 16, 0, 9, -31, 31, -29, -29, -8, -20, -4, 31, -21, 20, -14, -19, 4, -7, -14, -28, 27, -31, -8),
    (-6, 21, 4, 2, -2, 16, -21, 1, -21, 16, 20, 16, -41, -20, -3, -7, -14, -17, 5, -34, -7, 31, 63, -15, 13, 9, 44, -43, 0, 37, -29, -31, -12, 7, -7, -14, -6, 5, 43, -17, 25, -11, 0, -10, 18, -10, 52, -16, -19, 7, -12, 14, -8, -24, 31, 43, -1, 19, 20, 6, -9, -25, 13, -3, -2, -3, 9, 14, -7, -17, 32, 31, 16, 21, 22, -46, -8, 20, 6, -15, -10, 22, 8, 4, 27, -4, -15, -10, 9, -15, 18, 10, -21, 1, -2, 31, -3, -17, -37, -2, 12, 11, 0, 17, 5, -58, -18, -8, -43, -18, 4, -30, 14, -46, 13, 11, 5, -29, 33, -1, 21, -25, 30, -11, 17, 16, -9, 24, -16, -9, -27, 12, 11, 16, 2, -40, 27, -47, -3, 34, 24, -17, -2, -2, -17, 19, 26, 24, -23, 27, 16, 8, 14, -28, 3, -50, -36, -23, -15, -2, 23, -8, -6, 11, -6, 9, 23, -57, 7, 21, -4, -9, 19, 25, -9, 4, -43, -25, 6, -4, -7, -28, 21, 27, 29, -8, 1, -4, -5, -19, -19, -21, 14, -7, -15, 18, -15, 10, -13, 19, 1, -6, -9, 24, -31, -14, -12, 6, 35, -6, 6, -10, -23, -13, 13, 1, -16, 10, -49, -21, 15, -5, -7, 13, 9, -5, 23, 14, -26, -2, 45, -16, -47, 29, 1, 16, 1, 0, -29, -13, -15, -28, -1, 25, -19, 23, 1, -17, 14, 22, -12, -4, 5, 9, -5, -15, -2, -12, 7, -27, -29, 8, -3, -39, 23, 10, -10, -14, 10, -13, -20, -40, -20, -51, 7, -9, -9, -38, 9, 10, -31, -8, 6, 33, 5, -17, -8, -8, 20, -7, 23, -6, -2, 40, 31, 21, 5, 29, 21, -38, 10, -22, -29, -5, 8, -35, 30, 6, -24, 10, 16, 4, 12, 13, 38, 30, 22, -26, 4, 10, -32, -5, 3, -28, 14, -16, -30, 22, 27, 28, 34, 2, -5, -9, -6, -10, 9, 13, 20, -32, 18, 10, -2, 9, -8, 5, 14, -23, -7, -6, -13, -4, -6, 25, 15, -45, -6, 14, -24, -2, 9, 2, 16, -21, 25, -4, 0, -23, -15, -2, -8, -5, -24, -27, 1, 32, -9, 20, -17, 4, -16, -21, 1, -15, 5, 14, -21, 3, 14, 11, 7, -19, 18, 13, 33, -23, -18, -26, -4, -18, -18, -14, 15, -14, -20, 16, -11, -31, 3, 13, 31, 6, 18, 3, -5, 13, -32, -10, -9, -18, 0, -33, 27, -17, 33, 47, 14, -23, 27, 4, -18, 1, -3),
    (32, 17, -1, 4, 29, 6, 8, 3, 5, 14, 13, -18, -19, 11, 9, 10, 4, -4, 18, -5, -16, 5, -12, -3, 6, -31, -12, 20, -27, -20, -20, 30, -18, -8, -16, 3, -15, -32, -22, -18, 34, -20, -17, -17, -22, -1, -22, 18, 13, 10, -1, -9, -13, 24, 12, 7, -2, -5, 7, -15, -18, -48, 5, -14, 13, -13, 35, 15, -3, 9, -1, 9, -8, -37, 43, 2, -23, 9, -21, -2, -9, 19, 17, -13, 5, 11, 20, -12, -21, -45, -3, -29, -15, -2, 14, 15, -1, 24, 30, 38, -2, -1, -13, 21, -20, -4, 18, -14, -25, -9, 15, -13, 36, -8, 10, 2, -47, -23, 27, -5, 33, -46, -14, 47, -36, 17, 16, 30, -7, -4, -26, -13, 7, -30, 23, -22, 2, 5, 12, 12, 0, -14, 33, -13, 22, 11, 23, 65, 10, 6, -5, 19, -27, 10, -28, -38, -6, -26, -27, -1, 37, 8, 30, -11, -12, -20, 41, -19, 2, -14, -2, 1, -22, -31, -2, -43, -35, -4, -4, 14, -30, -7, 36, -26, -2, 2, -1, 7, -11, 14, -11, -4, 28, 8, -4, 75, 1, -8, -8, 18, -5, 12, -25, 4, 27, 10, 1, -24, 42, 39, -4, 27, -42, -3, 23, -52, 17, -31, 7, 6, -14, -3, -17, 6, -36, -44, -50, -2, -8, -22, 39, 3, -5, 39, 9, 7, 12, 25, 18, 0, 42, -14, 11, 47, -32, -7, -19, -2, 30, 20, -16, -17, 39, 14, -8, 13, 11, 33, -7, 27, -9, -3, -22, -18, 7, -9, -27, 8, -8, -14, -26, -30, -21, -43, -5, -33, -1, -24, 19, -1, -12, -16, 12, -8, -7, 28, 7, -10, -3, 17, 19, 24, -7, 29, -16, 22, -38, -2, -17, -12, 7, -25, 13, -4, 21, -9, 28, 6, -8, 26, 4, -31, -5, -8, 25, 15, 1, -4, 11, 22, -25, 13, 16, -8, -36, 22, 21, -13, 51, 36, -4, -23, -5, -9, -22, -6, 28, -12, 25, 28, -7, 28, -21, -10, -4, -8, -8, -26, 6, 24, -3, 14, -13, -6, 21, -5, 23, 1, 19, -33, -25, -17, 22, -16, -17, -29, 2, 19, -13, -6, -26, 12, -36, -26, 29, -4, 26, -7, 0, 22, -5, 17, 2, -16, 38, -8, 17, 41, 14, -18, -17, -13, -8, 21, 20, -36, 18, 6, 20, 17, 17, -4, -30, 28, 4, 3, 32, -26, 5, -11, 30, -28, 5, -12, 6, 32, -35, -18, -29, -24, 15, -34, 8, -12, 21, -1, 0, 24, 9, 23, -9, 41, 9),
    (-5, 1, 24, 12, -29, 1, 23, -46, 26, 26, -25, -43, -3, -3, -42, 14, 6, -20, 3, 2, -37, -16, 14, 6, -29, 1, -3, 26, 11, 5, 11, -14, -44, -3, -30, -4, -50, -21, 7, 26, 60, 41, 41, 6, 14, -11, 15, -18, 14, -8, 4, 25, -8, -2, 7, -17, 0, -1, -9, -19, 17, 12, 7, 0, 13, -3, 1, 25, -30, 21, 17, -30, -21, -12, 17, -11, -17, 13, -32, -10, -28, 0, -18, 25, -42, 1, 35, -14, -4, 18, -16, 32, -27, -3, -1, 11, -17, -25, -34, 18, 1, -8, -15, 37, -9, -12, -21, 25, -17, -19, -16, -36, 22, 49, 23, -34, 3, -18, 21, -6, 26, -19, -46, -19, -23, -24, -25, -5, -39, -28, 28, 15, -18, -36, 30, -45, -3, -29, -50, -18, -3, 0, -8, 20, -5, 13, -15, 32, 3, -9, -15, -25, 9, 33, -50, -15, 35, 14, -18, 26, -6, -16, 15, -8, -12, -7, -5, -15, -57, -11, 29, 32, 37, -3, -14, 5, 35, -5, 24, 14, -15, -14, 4, 32, 6, -9, 73, -10, -26, 5, -29, 9, -4, 33, -12, -17, 6, 0, 1, -17, 36, 8, 6, -20, 38, -13, -7, 38, -5, 38, -38, -5, -29, -18, 14, 22, -46, 7, 1, 11, 16, 3, -6, 7, -30, -43, 25, 37, -17, -15, 14, 37, 21, 16, 30, 31, 3, 15, -17, -19, -9, 22, 14, 1, 0, 18, 14, 0, -10, 34, 29, 8, 12, -18, 2, 10, -1, -6, 15, -21, 7, -7, -5, -21, 2, 0, -21, -29, 3, 14, 31, 15, 4, 9, -20, 32, -9, -18, 14, -2, 10, 10, -27, -2, -6, 0, 1, -7, -20, 2, -7, 17, 10, -9, -20, -10, -43, -20, -15, 27, 12, -13, 1, 2, -5, 32, 22, -1, -31, -30, 17, 24, -39, -34, -2, -10, -5, -15, 13, 5, 2, -28, 25, 24, -14, -13, -3, -28, -7, -18, 5, -33, 3, 4, 8, 2, -17, 11, -31, -42, 6, -21, 12, -12, -21, 8, 21, 29, -9, 1, 19, -21, 14, 15, 1, -7, -2, 12, 4, 32, 11, 1, 15, -1, 19, -14, -11, -5, -1, -11, -21, 9, -5, -1, -18, 25, -13, -21, -17, 2, -2, 21, -26, -26, -23, 22, -2, 15, -12, 0, -23, -15, -16, 12, -12, 4, -7, 10, 3, -5, -22, -21, 17, 4, 3, -1, 22, -19, -11, 19, 25, 39, 10, 10, -2, 23, 13, 4, -13, -8, -2, 16, -13, -15, 11, 30, -17, -13, 10, 37, 42, -21, 8),
    (-13, 10, 14, -23, 1, -6, -3, 5, 8, -8, 29, 6, -1, 18, -17, -21, 25, 20, 8, 1, 35, -27, -23, -32, -13, -13, 13, -2, 23, -21, 26, 23, -5, 12, -12, -23, -25, -7, 30, 17, -19, 30, -22, -30, 12, -23, -13, -11, -2, -43, -25, -22, 18, -10, 1, 1, -18, 5, 0, -19, 10, 21, -30, -9, -11, -18, 3, 0, -8, -17, -37, -14, -17, 58, 5, -10, 15, 1, 15, -2, 6, -40, -6, -2, -4, -13, 29, -21, 39, 53, -7, 16, 14, 36, -18, -4, 9, 4, -26, -4, -35, -7, -34, -22, -21, 19, -8, -13, 7, 22, 3, -3, -20, 10, -15, -20, 56, -21, -21, 10, -19, 12, -33, -39, 3, -18, -12, -11, -6, 3, -31, -5, 16, -42, -19, -13, 11, 7, 0, 39, 10, 42, -8, -7, 12, -16, -8, 37, -28, 20, 8, 6, 11, 30, 24, 14, -11, 22, -21, -7, -39, -21, -18, -20, -20, 5, -12, -17, 24, 11, 17, -26, -43, -33, 18, 16, -13, -5, -24, 27, -20, -12, 49, 13, 6, -7, -23, -1, 18, -11, -4, -41, -17, 3, 18, 16, -28, 42, -20, 3, -5, 29, -8, -9, 16, 38, -25, 4, -37, -55, -5, -38, -44, -4, -24, -33, 16, 22, -14, 15, -5, -63, -19, 15, -8, -49, -43, 28, -13, -4, 31, -18, 39, 1, 19, 36, 31, 14, -30, -56, -26, 35, -5, 24, 3, -9, 7, -7, -24, 35, -3, 0, 27, 26, 4, -28, -22, -30, 11, 28, 11, 0, -5, 13, -40, 18, -16, -27, -2, -9, -34, -14, 25, -19, -25, -5, -6, -12, 3, -11, 19, -6, -6, 24, 37, -1, 0, -6, 18, 21, 13, -23, -4, 33, -16, 17, -11, 6, -36, 32, -62, 5, -5, -20, 6, -20, 21, -32, 20, 17, 1, -22, 4, -6, -1, -18, 13, 8, 10, -3, -37, -20, -17, 24, -2, -6, 29, -11, 0, 15, 19, 5, 17, 17, -9, -1, 15, 15, 1, -13, -17, -3, 2, 21, -1, -5, -18, 17, 34, 9, 42, -23, 0, -4, 9, -9, 5, 9, -11, 21, -10, 30, -49, 10, -7, -8, -19, -38, -20, -1, 22, -2, -14, 15, -22, -9, 31, -16, -24, -6, 6, 32, 29, -14, -12, -20, 2, 22, -2, -26, 11, 11, 13, -27, -19, 6, 13, 5, 20, -27, 43, -1, -40, 12, 31, 5, -36, -35, -37, 19, -13, 14, -31, 3, -1, -9, -31, -10, 10, -3, -24, 17, -4, 24, -24, -6, 29, -23, 31, 33, 44, -32, 14),
    (6, 18, -12, -16, 23, 4, 6, 12, 4, -28, 20, -7, -38, -23, -19, 28, 5, -11, 21, -20, -39, 20, 20, 20, -3, -9, 11, -36, -24, 35, 8, 11, 25, 35, 7, -9, 26, -8, 4, 7, 18, -22, -22, -18, -10, -22, 11, -39, -32, 41, 14, 11, 12, -16, 13, 8, -5, 28, 26, -19, -36, 6, -10, -21, -2, -32, 0, -9, 9, -20, 1, -33, 11, -7, -9, -31, -34, 8, 33, 27, 4, 26, 10, 21, 21, -16, 0, 12, -22, -23, -9, 15, 16, -18, -10, -21, -8, 6, 40, 8, -25, 4, -3, 34, 11, 20, -4, 7, -34, 2, -1, -11, -17, -20, 20, 7, -2, -10, 2, -26, -24, 9, 27, 13, -25, 24, 26, -10, 12, -23, 4, 4, -24, 11, 15, -22, -24, -29, -23, 12, 14, 27, -15, -7, -11, 2, 32, 36, 17, 1, -11, 28, -22, 47, -39, -10, -10, -8, 17, 31, -1, 10, -11, -50, -37, 6, -4, -19, 2, 16, -9, 11, -32, 20, -9, 16, 5, -10, -17, 11, 13, -42, 34, -18, 0, 1, -17, 32, -19, 16, -51, -44, -24, 33, 46, -13, -23, 15, 18, 8, 23, 44, -13, 7, -34, -9, 26, 20, -20, -34, -23, -40, -21, -11, 33, 3, -42, 25, 4, 10, 6, -16, 9, 10, 14, -12, 5, -3, 7, -22, -24, 3, -48, 20, 16, 22, 16, -7, -6, -30, 0, 34, 20, -12, -7, 32, -5, -15, -24, 24, 5, -30, 5, -23, -23, -38, 16, -5, -32, 36, -11, -10, 0, 4, -43, -13, 12, 12, -29, 0, 26, 16, 14, -28, -3, 32, 0, -41, 0, -6, 27, 20, 34, 9, 2, -13, 19, 15, 13, 44, 7, 9, -1, -27, -1, 53, -1, 3, 15, 13, -48, -6, 4, 11, -18, 17, -12, -5, -8, -1, -20, -13, 25, -13, 1, -35, -17, 14, -14, 5, -13, -1, 19, 0, 5, -3, 0, 16, -14, 22, -15, -49, 2, -1, 25, -14, -8, 19, -6, 2, -4, -1, 0, 1, -35, -10, -28, -23, 14, -12, 26, 33, 21, 2, 14, 12, -19, 14, -12, -13, -35, 18, 24, -15, -1, 29, -48, -33, 9, 19, -14, 15, -22, -2, 7, -33, 25, 16, 17, 6, -10, -1, 37, -36, 7, 40, 21, 31, -18, -8, -30, -12, 5, 20, 15, 8, 9, -40, -30, 30, 2, 3, -18, -33, -16, -16, 3, 13, -27, -16, -4, -11, 14, -16, 27, -44, -15, -58, 22, 58, 5, -25, 17, 17, -10, -2, -5, -17, 26, 5, 4, -8, 19),
    (-24, -25, -11, -36, -7, -20, -18, -49, -4, -21, 16, 17, 17, 24, -33, 5, -11, 12, 8, 10, -60, 30, 5, 22, -66, -23, -15, -8, 35, 40, -4, -5, -16, -2, -7, -12, 1, 22, -26, 0, 16, -19, 16, -29, -38, -15, -21, -3, -8, -46, 24, 4, 23, -25, -24, 3, 0, 10, 19, 3, -16, -12, -11, 9, 25, 46, 18, -19, -26, -19, 43, 39, -32, 11, 27, -2, 31, 0, 4, -5, 13, 1, -18, 20, -52, 36, -8, -3, -13, 5, 45, 10, -14, -10, -7, -29, -9, 10, -2, -11, -7, 34, -15, -11, 6, -29, 20, -24, -4, 9, -24, 10, 35, 28, 25, -38, -29, -19, 32, -8, -30, -5, -20, -17, 15, 25, -5, -19, 1, 9, 1, -17, -35, 9, -18, -3, 21, -44, 48, -31, 9, 5, -22, 23, 3, -11, -2, -3, 12, 11, -17, -16, -1, 18, 1, 5, 28, 5, 5, -14, 7, -15, 12, -8, -1, 16, -8, 18, 7, -2, -24, -4, -3, 3, 25, 24, 28, -7, -34, -24, 20, -11, 6, 9, -32, -9, -13, 6, -24, -39, -24, -4, -7, 17, 2, 6, -19, 18, -7, 33, -2, 6, -8, -12, -17, -5, -9, -3, -14, 53, -31, -40, 4, -1, 24, -2, 21, -10, 15, -27, -16, 11, -4, -28, -20, -12, -42, -13, -20, 33, -16, -35, -32, 17, 5, 8, 0, 20, 32, -22, 1, -9, 21, 8, 0, 13, -5, 17, -25, 11, 7, -15, -24, -26, -16, -12, 5, 5, -7, -52, -22, -8, 32, 2, 9, 6, -23, -31, 0, -1, 11, -4, -22, 14, -30, 36, -33, -28, 15, -26, 21, 40, 58, -21, 2, -2, -11, -27, 2, -9, -8, -29, -1, 11, 14, -42, 28, -3, -19, 42, 13, 35, -14, -12, 27, -31, -4, 15, -18, -18, -1, 12, -4, -9, -1, -37, -34, 11, 0, -12, -19, 13, -8, 25, -35, -23, 4, -10, -1, -21, -7, -4, 11, 9, 22, 10, 2, 6, 2, 13, -14, 11, 30, 1, -12, -11, 34, 21, -16, 29, -23, -22, 24, -34, 22, -14, 12, 20, 33, -19, 38, 30, -19, -22, -45, 23, 16, -26, -23, 15, -2, -26, -25, 3, 28, -15, 25, -9, -12, -9, -18, -11, -13, -18, 44, 7, 13, 18, -25, 15, -18, 33, 6, 42, -3, 14, -27, -11, 24, -24, 25, 0, -17, 3, -16, -7, -2, -20, -6, 49, 21, -9, -22, -34, 33, -21, -20, -32, -20, 11, -17, 18, 18, -19, 3, 0, 15, 16, -1, 18, 13, -52, 9),
    (17, 18, 15, -17, 13, 13, 16, 14, 9, -22, 4, 25, -33, -31, 15, -3, 14, 12, -17, -6, 1, -9, 28, -34, -11, 17, 3, 3, -17, -6, 22, 36, 1, -24, -9, 0, -4, -16, 25, -31, 17, -16, 32, 26, 38, 15, -24, -30, 30, 0, -20, 4, -23, 25, 18, 14, 0, 26, -6, 18, -24, 13, -16, -9, -2, -18, -10, 1, 16, 0, 57, 7, -14, 51, 16, 5, -22, -13, -4, 24, 26, -13, -12, -49, -10, -18, -2, 19, 18, -6, 22, 6, 29, 14, -41, -42, -25, -9, 4, 32, 23, 20, 6, -22, 2, -3, -23, 16, -37, -35, 2, 11, -9, 7, -25, -10, -12, -4, 22, -26, 3, 8, -13, -44, 25, -19, -27, -4, -26, -22, -11, 17, 16, -35, 13, -36, 15, 43, -14, 8, 21, -6, 5, -20, 1, -32, 2, -32, -12, 13, 17, -10, 21, -27, -19, -6, -1, 20, -5, -31, -7, 5, 31, 30, 13, 9, 22, 41, -18, -7, 19, -3, -6, 4, -13, 22, 45, 17, 34, 7, 18, 39, -17, 9, -25, 20, 0, -49, 30, 20, -16, 8, -28, 35, 22, -1, 3, -29, 13, 32, -9, 2, -7, -14, 21, 30, -29, 14, 9, 10, 37, 13, 22, 29, -5, -5, -28, -2, -27, -6, 37, 35, -18, 8, -6, -7, -20, -27, -16, 0, 0, -16, -22, 16, -15, 1, 40, 8, 6, 5, 9, -3, -24, 23, -3, -5, 36, -11, 31, 45, -9, -7, 14, -2, 31, -13, 1, 35, -17, 13, -11, 16, 24, 5, -18, 8, 3, 10, 25, 35, 26, 10, 22, 10, 17, -17, -11, -12, 38, -11, -20, 20, -9, 7, -9, -26, 28, -19, 11, 8, -17, -5, 27, -25, 5, 47, 13, -21, -42, 27, -27, 33, 7, -18, -28, 26, 15, -3, -51, 9, -15, -10, -5, -15, 3, -38, -15, 4, -1, -6, 12, 24, -19, 7, -1, -18, 3, -18, -12, -13, -13, -2, -18, -4, -2, 4, 16, -25, -17, -9, -2, 10, 5, -1, -27, -28, -22, 9, -22, 18, -4, 13, -20, 14, -29, 10, 19, -24, 40, -15, -2, 12, 23, -41, 4, 8, 2, 19, 18, -35, -21, -26, 16, -24, 10, -18, -1, -16, 4, -60, -5, -38, 3, 32, -10, -32, 6, -29, -8, -4, -17, 17, -30, -13, 9, -17, -22, 21, 14, 6, 9, 21, 14, 10, -12, 16, -3, 3, 0, 11, -2, -12, 8, -38, -19, 39, -34, 17, -17, -6, 19, 34, 30, 0, 14, 1, 2, -35, 26, 2, -2, 12, -3),
    (-8, 7, 48, -24, -15, 10, 25, 39, -37, 14, -28, -2, 23, -19, 9, -42, 1, -12, -12, -22, -26, 30, -35, -28, 61, 16, -5, 25, 5, 1, -14, 20, -18, -8, -16, 8, 6, 27, 9, -24, -10, 11, -48, 25, -18, 14, -27, -19, 19, 0, 20, -7, -10, -9, 7, 7, -34, 33, -16, -6, 48, -28, 17, -18, -6, -23, 0, -10, 10, 8, -1, -7, 34, 32, -21, -12, 9, -14, -12, -22, -19, 10, -12, -9, -4, 12, -1, 4, 16, -6, -7, 8, 28, -32, -12, -25, 25, -15, -12, -14, 16, 9, -23, -22, -37, -6, 26, -32, 23, -3, 12, 10, 8, 33, -9, -13, 40, -2, -13, -1, 5, 20, -14, -24, -22, -29, -12, 14, -19, 23, 17, 5, -25, -37, 24, -19, 9, -9, -8, -22, 12, 30, 16, 28, 21, 20, 11, -35, -2, -13, 31, 30, 18, -24, -8, 8, 25, 18, -3, -2, 4, 8, -21, -9, 3, 17, 13, 2, 24, 33, 26, 12, -20, 31, -10, 2, 15, -1, 37, 9, 33, 23, -8, -18, -27, -12, 16, -16, 38, -6, -6, -35, -20, 17, -10, -31, 15, -10, -2, 34, -5, -10, -6, 1, 41, 3, 37, -24, -7, -5, 21, 4, 17, 32, -1, -16, -10, 31, 20, -9, -8, 21, 10, -22, -8, -38, 2, -20, -35, 38, -22, 22, -25, -22, 17, -11, -2, 9, -34, 23, -7, -21, -6, 18, 30, -15, 32, 13, -29, 4, -10, 28, 14, 12, 29, -27, 5, -9, 15, -4, 4, -6, -19, 17, 12, 23, 20, -16, 33, 14, -5, 22, -24, 11, -3, -30, 0, 12, 9, -18, -14, -21, 20, -6, -15, -4, 18, 8, -3, -13, -6, -1, 4, -16, 7, 23, -23, -10, -7, 7, 4, 21, -7, -11, 7, 12, 7, -19, 11, 26, -18, 18, -12, -19, 5, 14, 25, 7, 6, -17, 3, 16, 18, 27, 25, -14, -17, 32, -21, -7, 18, 25, 26, -7, 11, 0, -12, 24, -3, -3, 19, 14, 16, 13, 35, 40, -22, -1, 18, -17, -1, -13, -10, -2, -30, 7, -15, -15, 5, -11, 3, -23, -3, -21, -27, -20, -54, 3, 3, -16, 31, -18, 6, -13, -10, 8, 2, -43, -27, 1, 43, 28, -29, -4, 8, 30, 18, -10, -22, 14, 22, 19, 8, 21, -6, 4, -7, -5, -6, -38, -45, 14, 34, 14, 14, 5, 32, -6, 3, -28, -22, -5, -10, 4, -23, 0, 20, 22, 20, -15, -28, -14, 17, -7, -60, 19, 17, 0, -20, -12, -21, 18, -9),
    (-2, 42, -29, 20, 3, 15, -6, -20, -18, -18, -4, -21, -56, -27, 18, 13, -9, 1, 18, -22, -23, -30, 22, 20, 2, 26, -4, -31, -39, -34, -37, -36, -30, -9, 18, 1, 2, 17, -37, 3, 18, -19, 9, -16, 22, -33, 20, 45, 14, 35, -18, 31, 21, -19, 16, 10, -17, -5, 14, 13, -37, -22, 18, -8, -17, 12, 23, -19, -20, -8, 55, 25, 15, 9, 24, 7, -5, 17, 7, 21, -22, 27, -4, 7, 26, -4, 14, 3, 22, -15, 13, 29, 4, -8, 1, 15, -23, 45, -20, 8, 2, 7, -27, 33, 16, 31, 3, 11, -19, -12, 28, -34, 2, -16, 5, -35, 2, -7, -2, -18, 17, -18, -2, 21, -27, 15, 12, 6, -4, -4, -42, 16, -15, -19, 7, 4, -23, 22, -12, -24, -3, -38, 2, -38, -38, 7, -16, -24, -16, -21, 6, 37, 29, -19, 28, -15, -13, -5, 3, -22, 12, -18, 22, -12, -17, 7, -21, -2, 4, -40, 10, 5, -28, -2, 14, -1, 20, 11, 19, 21, 19, -11, 8, -7, -1, 38, 4, 0, 12, -4, 14, -38, 4, 43, 9, -1, 10, 14, -29, -3, 11, 10, 23, 43, -29, -40, 34, 6, -33, -3, -19, 2, -8, 6, 13, 6, -21, -16, 5, 10, 8, -3, 22, 6, -14, 5, 32, 17, 12, 22, 9, 23, -10, 7, -6, 8, 29, -31, 15, -28, 4, 36, 19, 6, -35, 8, 17, 52, -42, 5, 5, -3, -51, -15, 34, -49, 1, -31, 4, -36, 4, -9, 17, -33, 13, -26, 7, -6, -15, -12, 1, 25, 20, -2, -22, 30, -6, 7, -4, -16, -42, 3, -22, 4, 28, -38, 49, -30, 14, 25, -12, 20, 20, -19, 5, -6, -12, -8, -3, -16, -18, 8, -4, 35, -29, -22, -32, -22, 10, -15, -23, 19, 3, -2, 13, 0, 2, -2, -11, 11, 7, 18, 30, -14, 18, -3, -30, 6, -11, 8, -34, -19, 0, -26, 1, 2, 21, 6, -17, 43, 5, -19, -15, -1, -17, -37, 3, -1, -39, -27, 0, -32, -1, 22, -16, -11, 20, -33, 5, 16, -11, 21, -13, -26, -3, 16, 7, -39, -11, -29, -36, -39, -8, 4, 25, -9, -33, 5, 11, 5, -21, 7, 21, 7, 18, -7, -26, 43, 5, -16, 8, 23, 15, 15, 16, 11, 13, -30, -18, -37, 8, -2, 1, -25, -28, -4, 15, -10, 4, -3, 2, 23, -40, -27, -16, -26, 8, -21, -18, -10, 6, -25, 8, 4, -5, 15, 21, 23, -21, 9, 35, -8, 7),
    (5, -21, -13, -10, -12, 14, -20, -18, 19, 43, -1, -4, 27, 18, 6, 42, -14, 16, 36, -9, -34, -5, 40, 4, -15, -36, -2, -24, 30, 13, -2, -6, 27, 3, 18, 21, 8, 15, -29, -43, -29, -20, 59, 18, -28, 22, -36, -45, -23, 43, 26, -17, -16, 6, 23, -19, -12, 34, 22, 33, 31, 16, -6, -8, 11, -20, 2, 17, -8, -21, -17, 26, 21, -39, 26, 10, 21, 10, -7, 21, 12, 34, -28, -12, 2, 38, -56, 13, -15, -14, 18, 18, 0, -12, -9, -33, -1, -9, 13, -5, -6, 36, -15, -18, -3, 29, -19, -1, -20, 7, 9, -10, -12, 0, -8, 2, -12, -15, 14, 23, 3, -16, -6, -21, 4, -6, 18, 26, -19, -19, -40, 18, -27, -18, -11, -3, -36, -12, 7, -27, -4, -12, -13, 1, 3, -4, -4, -13, -4, -25, -22, 12, -40, -19, 32, 26, 4, 1, -13, -28, 8, 35, -22, -1, -31, -22, 32, -8, 34, -1, 3, 0, -23, -8, 15, -9, -26, 12, -6, -28, -13, 17, -13, -6, -4, -10, -8, -28, -25, -19, -11, 12, 4, -10, -51, 25, 1, -6, -24, 48, -7, -13, -7, 10, -9, 19, -26, -32, -34, -8, 12, -17, -50, -12, -7, 22, 47, 28, -20, -26, -18, 11, -20, -4, -25, 11, -23, 19, 12, -11, 13, -43, -8, -2, -25, -22, -5, 5, -36, 11, 3, 11, -30, 2, -5, -2, -2, 4, -13, -8, -10, 7, 0, 4, 35, 1, 1, 42, 0, -2, -23, 1, -9, -16, 38, -19, -12, 16, 1, 5, 29, -13, -21, -12, -24, 15, 0, -42, 2, -36, 3, 22, -12, 17, 4, 20, 6, 10, 29, 14, -18, -13, -4, 25, -21, 0, 2, -4, 17, 24, -16, -21, -9, -25, 15, 0, 30, 27, -17, 1, -1, -26, 11, 25, 35, 13, 4, -6, 31, 1, -12, -25, 34, -8, -7, 22, 17, 9, 2, 31, 20, -40, -12, -20, -4, 26, -25, -20, -8, 3, -7, -11, 19, -37, 25, -6, -7, 1, 20, 6, 8, -10, 32, 16, -31, 5, 0, -3, 2, -6, 1, 7, 2, -13, -23, -2, -8, 12, -4, -61, 10, -25, 40, 39, 3, 10, 29, -11, 2, 12, 29, -5, 30, -23, -31, -7, -4, -2, 7, 6, -5, 16, -20, -7, 9, -16, 19, -6, -23, 1, 8, 23, 19, -23, 2, -17, -45, -15, -5, -9, -7, 42, 10, -24, 9, 12, 19, 5, 32, 27, 13, -10, 15, 1, 19, 16, -26, 29, 27, 19, 10, 7, -1),
    (-32, -22, 19, -36, 27, -13, -9, 26, -4, -7, 5, 26, 30, 6, -13, -37, 34, -2, 41, -10, 3, -10, 14, 9, -12, -29, -20, -1, 29, 25, -28, -9, 7, -19, 14, 5, -52, -10, -37, 12, -15, -30, 36, -11, 9, -9, -16, -14, -16, -24, 7, -26, -11, -9, 17, 0, 30, -21, 4, 35, 29, -25, -9, -18, 40, -30, 5, 13, 9, 27, 18, 23, 26, -18, 25, 13, 15, -7, -26, -52, -20, -4, 31, 11, -9, 52, 19, 16, 9, -41, 16, 37, 11, -21, 7, 7, -14, 1, 11, 43, 7, 22, 28, 2, 25, -21, 8, -3, -5, -5, -7, 16, 12, -16, -27, 18, -30, 11, -27, -18, 11, -14, -22, 5, -22, 1, -8, -4, -37, -24, 20, -14, 28, -32, 21, 20, 10, -17, 2, 14, -51, -22, 45, 15, -11, -33, -7, -7, 15, 0, -20, 30, -19, -9, -45, 33, 2, 1, -12, -2, -3, -11, 14, 10, 13, 13, 14, 22, -15, 15, 12, 16, -14, -4, -40, -41, -6, 0, 33, 3, -38, 11, -8, -3, 11, -19, 25, -10, 6, 15, -23, 6, -16, -5, 21, -2, 16, -29, 8, 2, 17, -2, -25, 16, 20, -3, -24, 2, -3, -21, -10, 44, 10, 21, 15, 30, 12, -23, -22, 25, -15, -10, -37, -33, -20, -23, 3, -20, 6, 57, -28, 27, -13, -40, 22, 20, -18, -4, -9, 1, -8, 3, 7, -23, -11, 13, 33, 24, 10, -22, -8, 0, -11, -43, -28, -6, 6, 18, -9, -8, -11, -8, 3, -3, -3, -22, 29, 30, -20, -13, -12, 11, -37, 2, 13, -11, 0, 54, 7, 29, 26, -16, -1, -22, -26, -7, 14, -28, -2, -29, 13, 5, 19, 6, 20, 2, -6, -16, 12, 1, -6, 19, -16, 8, 19, -12, 18, 25, 12, 25, -3, 17, -24, 18, -4, 9, 11, -14, -18, -12, -22, -23, 5, 49, -21, 13, -7, 36, -2, -31, -8, 7, 7, 11, 15, 43, -11, 27, 35, -35, 9, -8, 27, -40, 19, 4, -12, -2, 34, -16, 9, 11, -3, -9, -3, 26, -17, 11, -10, 11, 5, 6, 7, 3, -25, -10, -22, -12, -6, -15, 6, -35, 4, 22, 30, 39, -18, -15, 13, 15, -15, 12, -4, -19, 41, -26, 38, -14, 21, 15, 30, -3, 18, -12, 21, -26, -17, -30, 10, 36, -40, 23, 12, 15, -27, -3, 4, 3, -17, -20, 32, 7, -23, -45, -19, 17, -16, -5, -7, 7, 34, 7, 17, 6, 0, -31, -9, 24, 8, -19, 27, 3, 6),
    (-19, -13, 1, -2, 12, 9, -23, -7, -4, 1, 5, 4, -5, -5, -25, -26, 32, 3, 13, 10, -45, 1, 15, -18, -14, 1, -2, 26, -4, -8, -10, -6, -21, 6, 4, 41, -23, -7, -21, -29, 19, -35, 11, 14, -28, -18, -11, -22, 3, 23, 4, -28, 18, 46, -14, -28, -16, 34, 2, -1, -4, 14, 5, 8, -8, -12, -23, 15, -4, -13, 33, 11, -37, -1, -14, 24, -9, 17, -13, -34, -2, -3, -10, -1, 8, -19, 13, -28, -35, -4, 13, 21, 13, -2, 9, -19, -20, 7, -5, -3, 4, -3, -36, 14, -28, -1, -1, -26, 34, 21, -13, 10, -1, 31, -18, 7, 24, 3, 10, -6, 46, 12, -4, -30, 1, 9, 0, -6, -8, 2, -3, 27, -12, 19, 8, -21, -32, 11, 8, 17, 11, -22, 7, 21, -2, -8, 19, -13, 8, -7, -14, -19, 24, -56, -37, 7, 17, -4, 6, -49, 47, 11, 35, 19, -14, 26, -21, 40, 20, -24, -35, 9, 14, -14, 0, -30, -41, 8, 36, -14, -35, 51, -13, -10, 24, -65, 16, -7, -44, 20, 27, 5, 30, -19, 21, -30, -8, 2, -12, -41, -14, -21, -53, 7, -14, 16, 26, -30, 12, -47, 32, 39, 15, -12, 30, 36, -17, -44, -46, -27, -5, 8, -15, -7, 16, 19, -28, 37, -49, 34, 27, -22, -26, 11, 14, 1, -37, 5, 35, 7, -7, -19, -16, 0, 28, -16, -29, -14, -18, -12, -17, -1, -7, 35, 7, -11, -6, -19, -17, -10, 4, 32, 39, 19, 6, -20, -15, -14, -8, -16, 16, -31, 12, 36, -7, 28, -9, -4, -39, -7, -7, 18, -15, -19, 3, 30, -21, 15, -28, 46, 10, 13, -17, 6, -19, 0, 12, 3, -45, -34, 21, -20, 6, 29, -15, 18, 4, 46, -44, -23, 6, 3, 23, 14, 29, 33, 36, -52, 5, -24, -4, 0, 3, 1, 5, -7, 32, 12, 11, -14, -5, -11, -33, -21, 32, 10, -38, 4, 31, 7, -4, -22, -7, 24, 38, 8, -29, -40, -17, -5, -22, 21, -31, 21, 0, -3, -27, -9, 5, -12, 14, 2, 25, 20, 19, -13, 6, -41, 22, -7, 3, -22, -37, 29, -25, 1, 16, -8, -30, -24, -27, -5, 9, -22, -21, 12, 32, 3, -53, -35, 21, -3, 8, 22, -21, 7, 39, 5, 15, -27, 24, -2, -17, -1, 22, -31, -5, 9, 7, -29, -30, 25, -33, -23, -5, 2, -7, 5, -24, 9, -48, 13, 4, -19, 20, 8, 30, -34, -33, 16, 12, 17, 10),
    (-5, -6, 24, -46, 13, 11, -21, 6, 11, -7, 2, -8, -19, -12, 12, 7, 10, -20, 7, 5, 13, -2, 57, -23, 23, 1, -6, -15, 12, 23, -2, 4, -23, -3, 4, 14, 23, 54, 12, 22, -28, -18, -23, -21, 16, -11, -37, -33, 5, 13, -2, 18, -21, 21, -16, -14, 2, -1, -7, 1, -4, -19, -14, -14, -6, -3, 5, 40, 10, 10, 44, 14, -8, -34, 36, -6, -20, 23, 7, 9, -16, -35, 19, 36, -11, 3, 11, -28, 8, -1, 17, -26, 38, 11, 14, -4, 23, 15, -7, -17, -13, 24, -20, -12, -13, -16, 9, 26, -2, -11, 9, 3, -19, -11, -4, 25, 39, -3, 35, 17, 6, 4, -17, -7, -20, 11, -6, -26, -16, 10, 1, -9, -10, 9, 12, -10, -44, -22, 7, -4, -17, -6, -1, -17, 21, -37, -21, -3, -22, -11, -9, -3, 17, -42, 20, 4, -14, 0, 32, -36, -18, -15, -5, 35, 3, 21, 13, -3, 16, -19, -7, 10, 10, 10, -26, 13, -12, -24, 26, 0, 30, 27, -28, 9, 18, -44, -19, -24, 11, -35, -9, 34, 23, -5, 3, -1, -5, 14, 24, 5, 22, -12, -42, 18, 17, -15, -9, -8, -8, 4, -2, -4, 0, -9, -15, 14, 3, -12, 15, 12, 35, -21, -57, 6, -22, -15, 0, -7, -18, -11, 7, 9, 21, 8, 31, 27, -16, 12, 14, -10, -19, -27, -11, 34, -6, 28, 5, 23, 22, -3, -17, 7, 18, -17, 7, 18, 22, 21, -19, 17, -11, 1, 37, -27, 21, -36, -27, -44, 40, 4, -3, -27, -53, -33, 23, -7, -10, 2, 37, -25, 3, 10, 22, 5, 1, -18, 21, -30, 7, 12, 30, -4, -21, -31, 39, -22, 8, 15, -20, 26, 5, 9, -4, -4, 4, -14, 15, -15, 9, 23, -1, -5, 14, -20, -8, 17, 16, -20, -11, 13, 0, -10, -34, -26, 24, 4, 12, -3, -29, -7, -3, 29, 13, 33, -29, 6, 11, -13, 8, -7, 1, -23, 22, -31, 30, 10, -17, -38, 11, 23, 23, 28, -19, -25, -10, 24, 34, -25, -9, -27, -37, -21, -12, 45, 12, -30, 26, -9, 17, -48, -33, 17, 12, 25, -44, 15, 20, 11, 26, -3, -19, 30, 21, 22, -35, 23, -15, -9, 1, 3, 12, -15, 21, 41, 19, -26, 8, -5, -26, 27, -27, -19, 14, 6, -13, -25, 14, -20, 3, -18, 23, 29, 19, -7, 3, 1, 4, -4, -20, -4, 6, 14, 6, 36, 21, -20, 10, 0, -15, 28, 25, -12, -14),
    (9, 11, -29, -17, 9, 10, 27, 37, 5, -15, 27, 28, -13, 32, 8, 31, -38, 9, -19, 25, -16, 22, 7, 7, -14, 3, -10, -16, 2, -10, 14, -1, -22, 28, 22, -27, 52, -34, -13, -11, -8, 11, -6, 15, 21, -15, -67, -19, 8, 26, -37, -17, -30, 18, -17, 3, 10, 41, 29, 23, -10, 4, -7, 11, 5, 1, 0, -13, 13, 4, 4, 0, -7, 46, -12, -31, -4, -35, -39, 14, -8, 15, 20, -4, 13, 14, -4, 24, -14, -22, 14, 22, 1, 14, 35, -3, -15, 9, 6, 1, -14, 13, 23, -34, -20, 4, -13, -9, 2, 24, 30, 31, 8, 17, -6, 13, -18, 26, 13, 8, 7, 27, -4, -6, 5, 18, -31, 23, 21, 14, -13, -10, -8, 24, -22, 31, 38, 5, -36, 11, 3, 2, -6, -31, 27, -17, 17, 30, -30, 17, 11, 20, -2, -46, -30, 26, -36, 0, -7, -28, 30, 9, -48, -30, -13, -31, 69, 34, 31, 1, 17, 3, -39, 8, -31, -3, 9, -3, -6, 16, 1, 7, 38, -9, 18, -16, 27, -15, 3, 8, 35, -51, -12, -26, 19, -23, 6, -11, -22, 27, -18, -10, 10, 11, 2, -24, -9, 5, -20, 20, -24, -7, 0, -15, 35, 12, 31, 10, 11, -11, -15, 21, 1, 10, 20, 22, 19, 10, 17, 7, 50, -16, -13, -45, -4, 39, 4, -7, 16, 21, -17, -8, 2, -11, -22, -22, 6, -27, -8, -4, 38, 20, 8, 14, 28, 0, -33, -6, 11, -8, 0, -17, -2, 20, 17, -22, 12, 22, 16, 17, -26, -15, -4, 14, 17, 20, -19, -1, -13, -12, -29, 4, -10, -6, -23, -19, 5, -13, 8, -17, 12, 31, -1, 36, 40, -14, 13, -11, 16, 5, 2, -25, -32, 32, 1, 2, -16, 14, -1, 2, 43, -46, -9, -30, -33, -44, 28, 8, 0, -15, -25, -1, 13, 27, 6, 30, -3, -5, -10, -35, 66, 22, -25, -27, -14, 12, 17, -1, 49, 33, 6, 11, -6, -30, 5, 34, -18, -30, -6, 6, 20, -13, 31, 24, 31, -33, -22, -12, 6, -8, -6, 19, -28, -10, 13, 29, 2, 26, 16, -5, -17, -2, -13, -25, 18, 28, -18, -16, 43, 24, -37, -29, 21, 7, -18, -14, -5, 21, -5, 7, 3, -19, 4, 25, -15, -39, -12, -13, -26, -6, -40, -15, -10, 5, -1, -32, 9, 9, 6, 8, -25, -15, -41, 11, 10, 21, 24, 10, 12, 18, -38, 9, 40, -14, -14, -2, -10, -6, 13, -6, 6, 7, -11),
    (-9, 10, 1, -4, -27, -29, 2, 20, 17, -2, -14, 26, -48, -11, 3, -12, -3, -11, -12, -4, 30, -9, 1, -45, 8, 1, 5, 0, -13, 32, -19, -4, -40, 4, -38, -10, 5, -48, 7, -11, -10, 2, -44, 20, 17, -8, -20, 2, 8, -21, -24, -34, -1, -28, 7, 2, -23, -22, -23, -38, 26, 36, -4, -11, 9, -25, 0, -10, 20, -12, -34, -6, 10, -15, -31, 19, -4, -19, 10, -24, -1, -30, -18, -16, -23, -12, -19, 16, 6, 45, -35, 20, 19, 14, -7, 12, -20, -11, -42, 21, -17, -9, -4, 0, -18, 4, 11, -25, 15, 5, -20, -19, 15, -3, -18, -8, 23, 20, -15, -26, -22, 36, -10, 4, 8, -13, -10, -13, -13, -31, -48, 3, 25, -33, 17, -31, 34, 6, -36, -18, 15, 25, -17, 31, -26, 31, -19, 2, -11, 15, -27, 31, -5, -17, -19, -9, -6, -17, -30, 13, -53, -24, -16, -42, -26, 20, -21, 5, 40, 2, -5, -1, -51, 6, -10, 37, -39, 5, -12, -39, 38, -38, -2, -33, 5, 40, -52, 36, 10, -50, 3, -26, -14, 37, 18, -5, 1, -4, 24, 35, 20, 2, -5, -24, 4, 30, 15, 21, 39, 11, 14, -6, -10, 9, -12, -5, 21, 17, -19, 12, -1, -17, -9, -6, -14, -30, -22, 16, 4, -52, -5, 18, -17, 35, -23, 26, 30, 13, -54, -4, 8, 5, -25, 8, -20, 21, -8, -29, 13, 21, 24, 15, 53, 37, -22, 0, 1, -31, -5, 32, 14, 21, -3, -23, -12, 25, 0, -17, -35, -43, -6, 20, 10, -7, 1, -18, 26, -38, 21, -27, 15, 53, -2, -16, 40, 7, 22, 7, 1, 1, -23, 23, -9, -39, -21, -9, 8, -3, 22, 37, 19, -3, 16, -18, 4, -9, 8, -41, -20, -16, -41, 22, 19, 7, -14, -26, -14, -2, 5, 9, -5, 0, 32, -7, -14, -4, 12, -56, 1, -12, -19, 18, -16, 2, 15, -13, 1, 4, 9, 22, 4, -37, -12, 31, 10, 4, 7, 18, -21, 38, 29, -25, 33, -20, 0, -22, 50, 0, -7, -14, -8, -25, -41, -28, -10, -13, 31, -30, -21, -15, -26, 15, -10, -12, 33, 4, -5, 28, -26, 20, 2, 25, 27, 13, -13, -10, -2, -22, -30, 28, -25, -11, 14, -1, 13, -10, 21, 42, -3, 18, 22, -36, -4, 2, 43, 12, 4, -40, -33, -13, -2, -18, -7, -25, 18, -1, 45, -14, -25, 16, 0, -34, -6, 0, -11, -9, -4, 40, 18, 25, 24, 20, 22),
    (-43, -2, -41, 1, -3, 1, 21, -21, 47, -5, 9, -24, 19, 13, 21, 1, -63, 0, 15, -9, 5, -16, -69, -10, 0, -35, 7, 18, 11, -16, -4, 15, 19, 6, -45, -9, 0, -25, -16, -27, -23, 26, -12, 20, 4, -9, -20, 7, -1, -33, -46, -18, 0, -42, -2, -33, 33, -9, 20, 8, -26, 29, -12, 26, -27, 22, -9, 14, 9, 8, -35, 20, -18, 19, 8, 29, 22, -35, 18, -3, 1, -12, 8, -6, 25, -15, 17, 10, -3, -13, -20, 34, -8, -14, 5, 12, -5, -36, -22, -31, -19, -34, 2, -22, 20, 9, -18, -3, -29, 7, 1, 3, -43, -15, 26, 29, -14, -11, -38, 20, 0, 5, -25, -6, -9, -8, -30, -10, 17, -39, 13, -6, 12, 8, -3, -25, -5, -21, -4, 6, 19, 12, -30, 51, -17, 22, -43, -2, 24, -12, 1, 3, 24, -42, -16, 14, -26, 28, 28, 19, -34, -20, 34, 28, -1, 26, -12, 39, -19, 7, 14, 18, 28, -53, 5, 25, 8, 41, 10, -15, -24, 10, 6, 0, -2, -22, 2, 13, -5, -9, 15, 12, -32, -14, 18, 31, 20, -35, 8, -7, -7, -40, -10, -5, 5, -26, -14, -21, 19, 35, -16, -12, 15, 22, -36, 14, -15, -13, 25, 12, 20, -36, 7, -10, -31, 1, -18, -33, 10, 4, -42, 7, 14, -13, 15, 18, 3, -16, 2, 0, 4, -29, 2, 21, -5, 13, -16, -27, 13, -23, 10, 10, -42, -11, -25, 33, 14, 27, -10, -3, 15, 16, -36, 14, -33, -6, 4, 10, 29, 16, 18, -23, -33, -17, 22, -9, 8, -20, 24, 27, 46, -6, 14, 17, -16, -6, 7, 31, -11, 14, -5, 5, 22, -30, 11, 6, -24, -15, -19, 22, 37, 37, 3, 6, 25, -20, 25, -36, -29, 8, -16, 25, 3, -34, 9, -21, -3, -16, 6, 1, -19, 1, -17, 18, -19, -20, -10, 11, -39, -55, 24, -20, 15, 1, -5, 9, 26, 26, 15, -19, -6, 10, 0, 16, -28, 8, 11, -6, 18, 0, -29, -16, -10, 10, 23, 0, -8, 11, -12, 12, -15, -14, -34, 5, 44, 1, -3, 11, 21, 7, -12, -8, 13, 29, 16, -31, -43, 9, -15, -3, -7, -14, 2, 35, -28, -41, -35, -12, -16, -2, -39, 5, 15, -3, -29, -37, -39, -12, 17, -8, -8, -11, 10, 19, -5, 12, -16, 0, -10, 12, -7, -3, 14, -15, 11, -14, 14, -3, 8, 32, -14, 29, 18, 16, -4, -23, 31, -11, 15, -17, -6, -12, 1),
    (-10, -32, 5, -26, -10, -33, -37, -16, -34, 0, -32, -17, 11, 34, 25, -34, 2, -22, -10, 18, -15, 14, 34, 31, 23, -26, 4, -16, 11, 1, 12, 9, 32, 18, 6, 10, -16, -26, 32, -22, 8, -10, 2, 2, 5, 0, 0, -26, 5, -34, -29, 42, -6, -7, -29, -1, -36, 7, 25, 13, 7, -1, -25, -19, 16, 32, -17, 6, 4, -7, 47, 4, 43, -13, 2, 26, -6, 11, -26, 16, 6, 15, 3, -15, -25, 7, -7, -25, -14, -22, 11, 11, -29, 0, 37, 8, -11, -8, -1, 45, -29, 1, -30, 8, -30, -23, 29, -18, -24, -34, 1, -1, 33, 1, 16, 23, -19, -32, 49, 11, 12, -15, -17, 11, -6, -12, -14, -4, 7, -15, 12, 13, -15, 15, 32, -19, 0, -30, 43, -12, -17, -27, 55, -4, 5, -1, -12, -8, -13, 4, -33, 2, -20, -33, -16, 11, 15, 13, -21, -51, 32, 7, 32, -10, 5, -9, 16, 23, -38, 21, -18, 6, -15, 39, -29, -26, -32, 4, 28, -21, -41, 34, 17, 37, -8, -58, 28, -26, -43, -13, -8, 12, 16, 3, 6, 7, -17, 15, -28, -2, 19, 15, -4, 17, 4, 6, -8, -22, 16, -22, 23, 8, -17, -15, 14, 2, -6, 9, 5, 5, -33, 20, 13, -9, -19, 14, -1, 19, -31, 27, 16, 2, 6, -28, 16, 11, -42, -5, 9, 21, 28, -26, -19, 40, 8, 23, 5, 15, -19, 14, -13, -28, -1, -30, -12, 9, -5, -18, -16, 23, 16, -22, 40, 0, 31, 30, 40, -20, -17, -16, -12, -32, 15, -2, -34, 23, 5, 5, -15, 6, 5, 5, 20, -12, -21, -23, 18, -1, -11, 35, 20, -20, 6, 13, 34, 38, 4, 26, 3, -10, 14, -33, 12, -4, -8, 27, 5, 12, -16, -24, 4, 9, 33, -1, 9, 18, 35, -22, -1, 26, -10, -14, -11, 4, 15, -19, 10, 9, -20, -2, -25, -17, -32, 4, 28, -25, -6, 23, 27, 6, -21, 24, -17, 36, -10, 3, 16, 21, 4, -2, 20, -29, 8, -6, 9, 9, 6, 16, -5, -32, 21, 12, 27, 33, -12, 5, -18, -28, 25, -19, 1, -23, -24, -15, 20, 2, 3, -26, -10, 9, -13, -19, -9, 9, -10, 9, 28, 32, -28, 4, -25, 41, -46, 11, 7, 33, -6, 33, -9, -1, -36, -41, -31, 4, -16, -3, -9, 13, 14, -14, 7, -25, -31, -20, -18, 5, -18, -14, 20, 15, -7, 28, 6, 19, 15, -4, 2, -5, -12, 21, -1, 18, 6),
    (-35, -10, -31, -39, -14, -9, 11, 12, 12, 8, -8, -26, -36, -25, -7, 47, 16, -22, -31, -7, -6, 19, -33, -5, -22, -8, 26, -17, -4, -19, -5, -14, -7, 54, 14, -7, 52, 11, -24, -30, 40, 15, -16, 7, -22, -51, 16, -33, -19, 32, -18, -75, 3, 7, 16, 11, -21, -4, -5, -2, -40, -12, 20, 45, -4, -2, -18, 14, 40, -23, -46, -25, -28, 28, -8, -19, -17, -4, -17, -13, -16, -12, 5, -14, 17, 5, -47, 8, 19, 25, 31, 1, -7, 4, -35, 37, -11, 41, -10, -38, -4, -21, -10, -17, 21, 24, 22, 11, -32, 35, 11, 7, 2, -21, -23, -6, 42, -6, -14, -10, -15, 6, -4, 14, 22, -6, -21, -29, 8, 17, 4, 1, -2, -17, 10, 9, 5, 35, 10, -6, 25, -2, -10, 21, -17, 20, -4, 43, 26, -39, 24, 63, -14, -18, -20, -10, -17, -12, 10, 33, 18, -7, 18, 8, -35, -15, 12, -9, 40, 16, -5, -36, -7, -6, 16, 1, -4, 27, 17, 0, 16, 33, -21, 14, 16, -13, 13, -41, -30, 1, 16, 6, 21, 27, 43, 24, 21, 4, 4, 37, -15, -36, -12, 2, -11, -44, 5, 45, 26, -18, 37, 2, 13, -10, 4, -16, 34, -13, 20, 10, -3, -16, -30, 11, -10, 8, -16, -2, -3, 33, -34, 10, 51, -24, 6, -16, 1, -45, 6, -3, -26, 10, 21, -7, -1, 17, -1, 42, -12, -22, -25, -4, -6, -23, -10, 24, 36, -33, 8, -7, 36, 11, 1, -9, -3, -16, 31, 22, -7, -29, -22, -23, -27, 37, -9, -26, -5, 18, 5, 0, 30, -10, -6, 12, -13, -37, -30, -5, 5, -4, 1, -1, 22, -3, -21, -27, 4, -12, -38, -26, 13, -3, -25, -12, -53, -12, -4, 41, -25, -4, 29, -20, -8, 15, -18, -10, -20, -3, 17, -20, 3, 8, 4, 6, -24, -30, -10, -18, 29, 14, -17, 10, 18, 28, -13, 39, 26, -35, -18, 16, 15, -4, -2, -28, -32, 24, 12, 24, 22, 15, -2, -24, -39, 37, -27, -22, 38, 3, 31, 14, 14, 13, -33, -12, -2, 12, 16, -3, -25, -33, 29, -25, -6, -4, -7, 9, -4, -29, -9, -9, 38, 12, 1, 50, 13, -14, -38, -3, -16, -24, -5, 4, 18, 9, -3, 4, 13, -24, -24, -12, -64, 16, 3, 10, 7, 3, -8, -2, 0, 31, 14, 6, -19, -14, -6, 9, -31, 9, -15, -21, 27, 10, -46, -1, 13, -8, 14, -4, 11, -23, -7, -8, -7),
    (-45, 38, 6, -33, -20, -6, -14, -27, -11, 4, 12, -20, -5, 40, -14, 21, -16, -35, 21, -19, -7, -8, 3, -3, -7, -23, -10, -38, -23, 17, 17, 2, 7, 24, -11, -14, -15, -34, -12, -1, 0, 49, 0, -15, -6, -30, -39, -13, -37, 50, 16, -30, -7, -42, -42, -11, 27, -1, 4, -7, 7, 29, -15, 24, -6, 29, 25, -4, 21, 3, 5, -13, -15, -25, -28, -4, -10, -28, 12, 4, 11, -8, 2, 10, 18, -23, -7, -39, -19, 28, -5, -22, -5, 13, -19, 5, 16, 34, 13, 10, 15, 19, 5, -22, -2, -8, -24, 11, -12, 16, 3, 18, 14, 38, -3, -31, 39, 18, -53, 3, -24, -4, -21, -2, -31, -29, 33, -39, -8, -8, 3, 12, 6, -26, -34, -5, 20, -4, 7, 4, 17, -11, -1, 0, -33, 17, -4, -11, 3, 17, 7, 19, 11, -10, -51, -17, 39, -1, -44, -13, 16, -35, 28, 12, -24, 19, -16, 21, 30, 16, -21, -2, -13, 0, -1, 18, 41, 4, -20, 4, 2, -55, -38, 13, 43, 30, -26, -4, -17, -26, -32, -20, -23, 30, 24, 29, 14, -12, -17, -35, -6, 23, -44, 5, 28, 12, 22, 16, 26, -6, -3, -11, -37, -3, -18, 13, 6, 32, -41, -5, -53, -36, -28, 25, 0, -24, 8, -4, -6, -28, -1, -31, -11, -8, -44, -37, -13, 7, -2, -8, 39, 28, -4, 25, 16, 9, 10, 24, -17, 26, 7, -13, -24, -29, -13, -2, 22, -5, -21, -20, 19, -26, -18, 15, 34, 6, -28, -26, -33, -17, 20, -7, 9, -8, -1, -12, -5, -25, 40, -22, -19, 17, -44, -12, -37, 22, 23, -22, -27, -11, 2, -31, -7, 16, -28, 6, 2, 20, -40, -40, 34, 27, -15, 16, 15, -10, 18, 37, -23, 6, -44, -1, -29, 22, -15, 21, -31, 2, -33, -13, 6, -20, 2, -1, -57, -29, -6, 9, 56, 15, 5, -45, 20, 45, 4, 3, 20, 34, -7, 9, 2, -19, -7, -22, -27, 24, -19, 19, 8, 3, -12, -12, 6, 21, -8, 41, 22, 7, 6, -11, -45, -8, 6, -1, -23, 19, -12, -34, -11, 11, -6, -5, -32, -28, 0, 16, 8, 4, -8, 5, 14, 49, 17, 36, 17, -14, 22, 4, -25, 9, -13, -35, -29, -34, 1, -1, -6, -22, -30, 5, 38, 19, 4, 30, 1, -18, -13, -42, -30, -3, -13, -3, -22, -9, 7, -5, 7, -17, 1, -4, -31, -7, 2, 6, 0, 29, 20, 26, 14, -1, 52, -40, 27),
    (-24, 21, -25, -38, -10, -30, -21, -48, 23, -18, -27, 15, -26, 24, 8, 1, -22, -14, 27, 13, -29, -4, -38, -12, 23, 2, 4, 11, 13, -5, -25, 16, 8, 4, -6, -14, -34, -17, -15, -36, -31, -20, -17, 7, -25, -7, 11, 2, -21, 26, 1, -58, 9, -32, -6, -1, 14, 1, -43, -11, -1, 11, 2, 2, 3, 2, 19, 10, 10, -2, -9, -4, -5, -17, -39, 35, 11, -26, -26, -10, 15, 33, -3, 37, -16, -20, -29, -33, 5, -11, -14, 10, 17, -6, 20, 13, 1, -5, -2, -47, 3, -12, -11, 9, 3, -27, -35, -33, 36, 24, 17, 9, 4, 6, -24, 11, 15, -19, -24, 25, -7, 6, -18, 15, 3, 6, -14, -10, 5, 29, 1, -2, -1, 0, -8, 35, -35, 16, 20, -41, -8, 39, -21, 48, -2, 19, -29, -28, 28, -21, 22, 20, -2, -36, 2, 17, 13, 25, 34, 44, -61, 28, 15, -22, -33, 3, -63, 49, 3, -53, 17, -25, -11, -10, 31, 22, -12, 37, 8, -13, -5, 11, -23, 26, -6, 30, -23, -25, -42, -10, -28, -3, -1, -25, -3, 3, 14, -44, -25, -7, 15, 29, 1, 1, -13, 18, 34, 4, 1, 6, 3, 30, 22, -10, -15, 13, 22, -34, 7, 18, -39, -19, 14, -5, 10, 11, -32, 1, 3, -8, -16, -38, -40, 16, 4, -47, -14, 31, -43, -22, -21, 7, 22, -9, 0, -6, 29, -4, -7, 1, 12, -2, -2, 22, -13, 14, -6, -14, -25, -13, 10, -35, -13, -15, 27, 11, -12, -20, 6, 21, -9, -12, 5, 9, -37, -10, 16, -25, 15, -53, -7, -2, -8, -17, 43, -22, 2, -5, -15, 6, -17, 14, 10, -19, 17, 28, 27, 10, -13, -11, 23, -2, -18, 14, -13, 5, 10, -52, -7, 4, -49, -32, 28, 1, 19, 22, -3, -2, -10, -15, 11, 5, -30, -34, 39, 9, -30, -20, -10, 18, -20, 15, -4, -41, -2, 14, 14, 7, -20, -33, -1, -20, 6, 6, 15, -2, 7, -14, 26, 17, 14, 15, -12, 1, -24, 22, 28, 12, -38, 14, -1, 22, 0, -22, 5, -51, 12, 18, -10, 7, -16, -4, -16, -32, -10, -1, -21, -14, -27, -17, -3, 22, -15, 11, 13, 4, 25, -9, 24, -29, -14, -8, -16, 30, 28, 0, -5, 0, 7, 18, 13, 7, -30, 34, 7, -19, -36, -22, 24, 22, -6, -20, -54, -33, 2, 10, -14, 0, 0, -3, 30, -53, 28, 44, -12, -17, 19, 6, 29, 21, 20, -9, 3),
    (-4, -21, 8, -10, 24, -39, 8, 15, -16, -45, 3, 31, -13, -7, -10, -13, 37, 7, 23, 12, -20, 25, 12, 12, -21, 5, 3, -3, -19, 23, 2, -11, 34, -14, 21, -19, 17, 4, -34, 21, -16, 18, -8, -14, 24, -3, 3, 30, -12, 0, -25, -10, -28, -27, 3, -8, 12, -59, -3, 7, -23, 14, -24, -29, 42, 24, -28, 31, -4, -23, -6, 25, -18, -24, 4, 9, 6, -17, 2, 12, -6, -16, 13, 9, 5, -23, 3, 4, -23, 24, -36, -34, -23, -31, -42, 43, 1, -18, -17, -7, 13, 20, -25, -33, -3, 11, 33, -18, -14, -16, -36, 5, 32, 11, -47, 3, -3, -22, -24, -2, 10, -29, 10, -9, -19, 20, 13, -21, -22, -48, -5, 27, 5, 15, 9, -12, -18, 26, 13, -16, -25, -5, -13, -26, 1, -6, 31, 24, 5, -24, -14, -2, -12, -23, -37, 3, -2, -11, -23, -27, -17, -20, 30, 20, 44, 1, -11, -18, 40, 23, -6, -1, -27, 24, -50, 22, -6, 1, 20, 15, 8, 34, 16, -23, -9, -24, -26, -14, 18, -23, -35, 45, 14, -12, 15, 20, -6, 21, 37, -10, 7, 15, -30, 48, -2, -18, -18, -31, 10, -2, 18, -35, 1, 33, 18, 11, 37, 28, 22, 26, -33, 27, -12, -9, -12, -14, -9, 2, 0, 43, 27, -8, -1, -27, 11, -12, 2, -19, 18, 8, -5, 24, 18, 31, 4, -14, 2, 23, 9, 6, -16, -6, -8, -27, -9, 4, 6, 22, -4, -3, -38, 6, 30, 0, 4, -2, 13, -33, -17, 0, 2, -10, -32, -25, -16, 12, -10, -18, -9, 14, 3, -51, -5, 17, 13, -23, -15, -1, 40, -18, 2, -7, 8, -23, 18, 24, -2, -7, -12, 28, -2, 3, 10, -23, 24, -45, 0, -10, 28, -15, -6, 22, 14, 2, -28, 19, -21, 2, 14, -17, 18, -24, 25, -30, -6, 29, 22, 11, -1, -13, -18, 27, 2, -25, -32, -14, 16, 15, 13, -10, -4, 16, 10, 20, -22, -11, 16, 43, -11, 9, 11, 5, -32, -17, 9, 5, 12, 24, 12, -23, -16, 31, -13, -2, 24, -12, -50, 29, -1, -6, 34, 13, -9, 21, -32, 2, -17, -18, 11, 13, -2, -28, -24, -12, -35, 29, 2, -5, -3, -35, 23, 25, -30, 26, -15, -3, 14, -15, 5, -26, 12, -28, 18, -21, -24, 4, -5, 15, 2, -4, -24, -25, -3, 11, -15, -34, -4, 18, 7, -21, -26, -7, -38, -16, -13, -30, 1, -14, -19, 16, -39, -5, -5),
    (-45, -13, -36, -32, -7, 8, 9, 16, 23, -36, -32, -16, -40, -21, 19, 18, 18, -27, -3, 33, -35, 5, -64, 17, 28, -34, 33, -7, -9, 22, -16, -20, -19, 35, 5, 12, 20, 12, 27, -1, 25, 18, -18, -7, -39, -48, -9, 44, -17, 3, -30, -5, -15, -22, 19, 13, 22, 0, -25, 32, 20, -2, -13, -13, -7, -39, 19, -38, -31, -7, -20, -28, 43, 15, 6, 28, -27, -9, -33, -37, -26, 6, -1, 1, -2, 31, 16, -36, -10, -51, -21, -7, -21, 7, -26, 0, -7, -29, -3, -43, -18, -39, -2, -25, -20, -32, -3, 25, -24, 8, -18, 0, -1, -17, 12, 6, 20, -11, -43, 20, -11, -35, 16, -22, -13, 13, -1, -2, -19, -5, 22, -6, 22, -3, -13, 18, 42, -10, -16, -19, 5, 12, 14, -8, -27, 33, -12, 25, -31, 19, -10, -10, 21, 9, 7, -3, -3, 6, 6, 34, -33, -3, 4, 11, 0, -1, -27, 1, -7, 9, 8, 41, 23, -31, 7, 24, 10, 16, -33, -20, 36, 10, -48, 17, 15, 13, 41, 19, -9, -25, -10, -16, -2, 43, -28, 23, 17, 16, 6, -2, 32, 8, 20, -24, -5, -10, 39, 27, -15, -24, -30, 4, -31, -2, -36, -8, 0, -20, 12, 26, 28, -18, 22, 14, 12, 18, -31, -14, 25, 17, -3, 18, -15, 17, -12, 2, 6, 4, 10, -11, 24, 3, -4, -1, -23, -40, 8, 19, -15, 4, -9, 24, 18, -22, -26, 14, 5, -22, -28, 4, 2, -2, -37, 12, 14, 15, -2, 7, -14, -12, -28, -28, 12, 33, -19, 20, 28, 28, 44, 19, 14, -10, -11, 12, 19, 21, -11, -17, -20, 12, -34, 9, -9, -27, -27, 6, -12, -16, -13, -13, 1, -19, 4, 28, -15, 20, -15, -7, -16, 17, -8, 11, -8, 23, -31, 14, 20, -26, 2, 12, -20, 34, -36, -26, -15, -41, 4, 13, 20, 15, 25, -50, 39, 0, 18, -9, 1, 36, -36, -15, 12, -3, 32, 39, -8, -8, 15, 24, 6, 1, -4, 17, -5, -25, -7, -9, -8, 7, 36, 11, -6, -12, 6, -2, 14, -11, 15, -10, -20, -22, -16, -37, -3, -13, 0, 22, 27, -24, 22, -15, 32, 29, 19, -26, -19, 26, -46, 24, -13, 12, -21, -14, -7, -4, 18, -34, -28, 18, -4, 2, 1, -3, 17, 6, -15, -18, -29, -7, 24, -22, 16, -28, -26, 2, 20, -16, -16, 14, 24, -38, -13, -19, 17, -18, 8, 42, 12, 12, 10, -35, 14, -13, -4),
    (-5, -24, -27, -54, -23, 15, 7, -45, -14, -8, 19, -10, -21, 41, 6, 41, -76, -32, 7, -2, -13, -2, -68, 24, -49, -18, -31, -15, -15, -13, 24, -19, 20, 5, 39, 18, -21, 0, 16, -15, 34, 27, -11, 17, 1, 18, -14, -1, 19, -31, 13, 11, 9, 17, -37, -35, 4, -19, 26, 15, -2, -2, 6, -37, 62, 26, -8, 7, 24, 36, 3, -14, -6, -6, -25, -26, 4, 17, -27, -28, 0, 16, -9, 13, -15, 31, -21, -15, -39, -17, -15, 8, -6, 3, 26, 33, 19, -11, 21, 22, 11, -14, -1, -34, -22, 3, -27, -36, 0, -37, -41, -7, 13, 28, -16, -27, -15, -1, 20, -27, -30, -27, 25, 16, -36, 11, 16, -21, 15, -11, -8, -22, -17, -37, -7, -7, -12, -26, 7, -1, -4, 19, 33, -27, 11, -13, -55, -23, -13, -18, 8, -59, -14, -4, -11, -1, 19, 37, -13, 39, -10, -31, 4, 34, 20, 36, -55, 9, -83, 3, -4, 2, 9, -44, 2, -56, -10, -14, 28, -6, -14, -6, -12, -15, 2, 27, -8, 11, 7, -11, 26, 10, 8, 10, -13, 21, -9, -46, -9, -68, 10, -5, 6, -1, 7, -6, 25, 21, 37, 1, -7, -13, 48, 36, 13, -5, -67, -49, 15, -3, -5, 5, 14, 27, -5, 2, -13, -31, -37, 19, 17, 13, -25, 2, 25, 9, -10, 25, 11, -14, -5, 29, 20, -17, 8, 0, -21, 4, -16, 0, -10, -25, 2, 18, -6, -2, 8, 26, -5, 3, 10, 9, -2, -26, -39, -1, 14, -14, 29, 14, -35, 7, 7, 13, -10, 26, -4, -22, -8, -7, -8, 22, 33, -19, -26, 15, 23, -3, 7, 5, 16, 2, -26, 2, -5, -5, 10, -8, -6, -20, 24, -16, -24, 16, -6, 21, -31, 6, -1, -17, -7, 9, -61, 11, 21, 1, 14, -2, -16, -17, 10, 31, 10, -15, -43, 8, 22, -5, 13, -26, 4, -14, -25, 20, 55, 29, -11, 15, 10, 10, 19, -33, -9, -4, -39, -24, 2, -4, 8, 13, -26, -3, 3, 35, -11, -31, 30, -28, -2, 11, 13, 17, -35, 1, -8, 15, 13, 13, -7, 18, -24, 1, -39, 0, 30, 22, -19, 7, 21, -38, -44, 22, 14, -15, -11, 35, 9, 26, 14, 19, -25, -2, -20, -16, -22, -26, 1, -35, -1, 3, 19, 15, 13, -15, 10, -32, 12, 18, 32, -21, 15, -16, 13, 17, 33, -11, 27, 28, -27, -11, -25, 5, -1, -57, -15, 17, -2, -47, -17, -14, 26, 3, 20),
    (-10, -34, -23, 11, -29, -20, -39, -3, 0, 9, -3, -19, 14, 15, 7, -23, 15, -15, 6, 6, -26, -10, -1, 2, -25, 0, -9, 21, -13, 0, -8, 32, -20, -13, -14, -26, 2, 0, -12, -4, 8, 20, -22, -3, -24, 3, -15, 31, 4, -7, 9, 12, -14, 5, -30, 10, 36, -12, -1, -1, -26, -3, 17, -16, 10, 15, -42, 9, -26, -53, -29, -8, -7, -20, 21, 10, -5, -22, 2, -6, -16, -8, 0, -11, 11, -16, -22, 24, -12, 9, -9, -3, -23, -6, 24, 18, -7, -26, -19, 19, -6, 14, 2, 15, 1, 30, 23, -22, -6, 11, -9, 9, -30, 28, -28, -13, 4, -41, -15, -61, 7, 0, 2, -4, -32, -27, 21, 9, 17, -15, -35, 17, -11, -22, -5, -28, -34, 25, -10, 20, -2, 7, 17, -7, -19, -1, 15, -23, 13, 4, -19, -11, 5, 24, 21, -29, 27, 27, 11, 48, -30, -12, -1, -27, -1, 5, -27, 16, -25, -15, 2, -3, 37, -12, -19, 23, 24, 9, 5, -32, -19, 20, -44, -27, -1, -39, 11, -8, -4, 9, -19, 19, -43, 32, -19, -30, -16, -12, 31, 0, 22, -9, 9, -28, 2, 3, 6, 44, -36, 4, 8, -7, 38, -5, 1, 18, -28, -11, 37, -15, 34, 28, 34, -27, 37, 12, -5, -2, -3, 23, -11, -5, 41, 30, 47, -2, 12, 35, -12, -8, -5, 14, -56, 6, -11, 4, 34, 21, -4, 11, 23, -22, -12, -15, 18, 27, -7, -15, -27, 11, 12, 19, -36, -21, 13, 33, 17, 1, 3, -2, 6, 10, -13, -20, -1, 2, 23, 29, 2, -32, 43, 2, 14, -3, -10, -7, 11, -22, -16, 36, -24, 3, 2, -16, -20, -4, -16, 7, -8, 16, -16, -45, -17, 6, 21, -12, -23, 7, 4, -22, 32, 38, 31, 0, -13, 18, 7, -3, -18, -29, -17, 14, 10, 13, -5, -14, 13, -10, -12, -13, -7, 3, -33, -48, 12, -10, 15, -23, 6, 18, 10, 5, 11, 25, 17, -11, 20, -26, -9, -4, 17, 7, -4, -6, 30, -11, -2, -22, 33, -3, 5, -8, -18, -39, 7, -8, 26, 28, -1, -4, -28, -16, 21, -18, 27, -10, 26, 34, 21, -2, 3, -23, 24, 10, -41, 6, -40, 35, 3, 35, -5, 10, -6, -29, -9, 0, 1, -25, -4, -17, -19, -36, -2, -15, -21, 9, 33, -16, -8, 9, -5, 13, -1, -32, 19, 15, -2, 17, -37, -28, -5, 2, 5, -15, 35, 17, 22, 10, 5, 0, -2, -1, -4),
    (9, -31, 38, -4, 40, 4, 15, 16, 20, 20, -9, 21, -7, 1, 26, 1, 7, -44, -14, -23, 10, 42, 25, -17, -26, 17, -30, -20, -4, -9, 3, -32, -10, 8, 11, 11, -37, -16, -12, -15, -52, -11, 27, 7, -31, -28, -21, -41, -11, 6, 17, -3, 13, -31, 31, -16, 20, 10, 1, 41, 24, 27, 36, 1, -11, -58, -5, -14, -1, 11, -14, 22, -7, 18, -11, -24, 17, 10, -19, -12, 13, 2, 28, 16, -30, 20, -11, -11, -1, -37, 60, 16, -7, -16, -30, -14, -7, -10, 9, 7, 14, -26, -5, 12, -14, -15, -33, 17, 27, 0, 2, -37, 13, -32, -3, -31, 28, 22, -39, 15, -22, 9, -20, 2, 3, 9, -8, 8, -24, 7, 22, -11, -18, 18, 14, -6, 1, -25, -25, 11, -2, -9, 2, 16, -20, -12, -26, 18, -25, 12, -31, 25, 10, -36, 1, -3, 35, 12, 10, -4, -18, 2, 1, -26, 21, 27, 19, 28, -25, 3, 23, -22, -7, -21, -17, -20, 16, 36, 9, -15, 11, 40, 21, -21, 10, -9, 16, -32, 18, 33, -14, 12, -38, 30, -16, 39, -18, 0, -12, -13, -4, -37, 19, 4, 7, 6, -13, 32, -59, 26, -17, 11, -24, 4, -18, 29, -10, -22, -10, 5, -19, -17, -5, 0, 12, 4, 7, 16, 16, 26, 9, 3, 10, 27, -26, -14, -18, 7, -17, 12, -17, 11, -6, 7, 4, 25, -9, 19, 1, 11, -19, -6, 12, 16, -14, 16, 26, 24, -9, -40, -23, -9, -35, 14, 16, -32, 23, 0, -16, 1, -16, 2, -6, -20, -1, 18, -15, -18, 36, -18, 5, 20, -26, -36, -7, 22, -15, 4, -12, -23, -26, 38, 16, -21, -39, 14, -14, -2, -9, -28, 35, -15, -1, 25, 0, -10, 3, 6, -4, -33, -28, -15, -8, -10, -1, 35, -12, 2, 42, -28, 25, -44, -14, 32, -1, -41, 0, 9, 2, 4, -14, 7, -3, 37, -6, 47, 30, -1, -20, 11, 14, -22, 8, -5, -9, -35, 25, 19, -27, -11, 13, 20, -3, 0, -12, -4, -31, 0, 12, -12, -22, 3, -11, -4, -6, -7, 30, -1, -12, -10, 1, 21, 3, -14, -38, -23, 22, -43, -1, -14, -24, -8, 14, -32, -3, 7, -16, -36, -20, -21, -29, 41, 18, 11, 15, -7, 1, -1, 12, -29, 18, 32, -28, -42, 25, 16, 18, 5, -2, 20, 14, -22, -17, -23, -26, 27, -29, -17, 3, -5, 38, -5, 0, 4, -10, 3, 11, 5, 0, -4, 1, -38, -2),
    (-5, -22, -11, 2, 20, -23, -35, 3, 0, -25, -25, -7, 26, 21, 19, -14, -6, -15, 13, -19, -24, 1, -41, -14, -2, -35, -13, 10, 21, -31, 17, -12, 41, 12, -17, 9, 38, -6, -18, -14, -3, -19, 18, 25, -60, 4, -5, 6, -22, 17, -24, -37, 13, 0, 15, -11, 15, -38, 9, 6, -26, 11, -19, -6, -31, -4, 2, 40, 8, 24, -1, 12, -17, 19, -7, 36, 26, 2, -7, -1, 17, 25, 31, 20, 27, 20, -16, 3, 29, -24, 8, 1, 12, -4, -22, 45, -27, 28, -40, -21, 0, 3, -16, 25, 18, -34, -14, -12, -37, -16, -2, -13, 0, 15, 14, 12, 0, 27, -17, 4, 10, 2, 27, -14, 6, 13, -19, -29, -4, 7, 21, -8, 26, 23, -2, 7, 4, -36, -20, 24, 12, -3, 31, 20, -26, 11, -13, -12, 26, -31, -38, 15, 27, -17, 12, 8, 6, -22, 25, -1, -15, -7, 0, -12, -12, 21, -16, 58, -10, 5, -33, 14, -12, 1, 0, 9, 11, 31, -3, -9, 30, 36, -11, -36, -31, -13, 2, -11, 3, -28, 2, 4, -10, -8, -20, -6, -28, -3, -3, 0, 27, -33, 32, 28, -15, -20, 12, -41, 11, 7, 30, 2, 5, 0, 13, 16, -1, 4, -21, -9, 13, -6, -32, -17, 0, -36, 14, 6, 22, 15, -2, 9, -43, -20, 1, -4, -25, 18, 25, 14, -22, 7, 11, 15, -1, -4, -29, -17, 15, 29, -26, 33, -11, -24, -6, -45, -24, 5, -37, -38, 7, 3, 41, 31, 14, -11, 21, 8, -17, 17, -5, -1, -29, -46, 12, 12, -19, -14, 36, 10, -45, -29, 16, -21, -10, -4, 11, -14, -26, 25, 20, 13, -31, -39, -6, 46, -4, 11, -21, 15, 18, 14, -23, 19, -13, 37, 10, -43, -7, -19, 22, 0, 20, 10, -16, 16, -23, -11, -7, 7, 6, -17, -28, -17, -16, 7, 26, 20, -53, 9, -28, -5, -26, -27, -22, -7, -7, 14, 5, 22, -27, -16, 25, 39, 38, -5, -10, -13, 11, 8, 7, 2, 7, -32, 15, -27, -19, -30, 22, -19, 9, -11, -22, -17, 20, -3, -2, 12, 5, -27, 10, 22, 16, -47, 26, 22, 8, -11, -1, 11, 32, -15, -20, 7, -7, -8, 16, 4, 22, 31, -2, 3, 35, 36, -34, 1, -6, 14, 37, 34, -30, -16, -21, -10, 26, 6, -9, -43, 22, -19, 17, 20, 16, -21, 14, -33, -21, -21, 33, -42, 21, 15, -5, -2, 5, 15, -27, 29, 14, -9, -8, -41, -9),
    (10, 15, 4, 51, -32, -8, -35, 4, -24, 31, -41, -14, -22, -29, 34, -17, 15, -23, 19, -17, -61, 9, -13, -17, 27, -11, -10, 22, -8, -8, -48, 7, -20, -33, -21, 23, -27, 20, -20, -21, 7, -3, -3, 1, -8, 2, 13, 13, 7, 4, 22, 0, -8, 46, -4, -2, 28, 35, -28, 49, 10, -9, -10, -45, 1, -29, 20, -31, -4, 4, -5, 36, -11, 10, 3, 15, -14, -25, -24, -9, 3, -2, 11, -3, 8, -1, -12, 16, -30, -21, 3, 15, -7, 0, 26, 52, -6, -18, -11, 21, 25, 17, -30, 18, -34, 38, -7, 26, 43, -52, 23, -16, 43, 52, -48, 7, -27, 41, 3, -37, 5, 19, -11, 31, 1, -19, -3, -33, -33, -63, -46, 29, -41, 25, 7, 21, -13, 26, 47, 24, -3, 33, -2, 3, -23, 9, 24, 45, -12, 20, -14, 11, -29, 38, -8, 2, 13, -13, 8, -19, -11, -6, -21, -32, -65, -5, 21, -33, -48, -28, -12, -14, 8, -13, 21, 2, -13, -32, -39, 0, -4, -19, 25, 8, -54, 20, 38, 17, -30, -14, 36, -17, -9, 4, 11, -23, -1, 37, 24, -20, 22, -10, -19, 13, 16, 9, -11, 3, -9, -32, 18, -34, 29, -16, -15, -1, -16, 22, -28, -32, -24, 24, 15, 0, -14, -36, -1, 17, 7, -27, -14, 4, -4, 7, 6, 26, -7, 6, 1, -28, -22, -13, 29, 29, -49, 35, 15, -22, 9, 31, 20, -14, 36, -2, -19, 23, -5, -33, -24, -1, 22, -2, 26, -10, -15, -12, 31, -37, 1, -15, -1, -4, 5, -25, -18, 20, 27, 1, 34, -30, 19, -10, 24, 30, -24, 14, 14, -7, 6, -8, -18, 9, -26, 22, -5, 9, -29, -23, -18, 18, -4, 6, 19, 0, -7, -17, 8, 18, 8, 27, 0, 0, -15, 24, 12, 15, -42, -8, 28, 19, 13, -9, 5, 5, 23, 8, 56, -3, -26, 15, 8, -26, 16, 22, 19, -39, 23, 9, 16, 24, 6, 12, 14, 6, 1, 25, 20, 34, 22, 32, -11, -22, -7, -29, -21, 7, -3, 3, -23, 15, -23, 19, -13, 1, -16, 0, -17, -15, -4, -15, 5, 22, -23, -7, 12, -6, -3, -5, -3, 16, 22, -8, 20, -40, -3, -52, 2, -16, -37, 0, -19, 21, 16, -40, 13, 18, 7, 12, 12, -31, 29, -4, 10, -7, -13, 7, 10, -14, -28, 14, -22, -16, 14, 22, -5, -27, 13, -14, 28, 4, -47, -11, -2, 29, 9, 7, 37, -18, 29, 21, 19, -20, 11),
    (-4, 30, -11, -19, -20, 8, -33, -8, 12, -9, 9, -14, -23, -6, -6, 30, 25, 0, -26, 4, -12, 14, 7, 8, 5, 16, -8, 4, -2, 9, -16, 1, 0, -18, -19, -17, -24, -52, -5, -21, 37, 55, -10, -21, 19, -7, -31, -1, -25, 56, -19, -21, -13, 22, -45, 2, -18, 16, 10, 3, 10, -9, -37, 1, 3, 17, -29, 30, -10, 20, 32, 24, -13, -20, -47, -44, 12, -2, -27, -16, 23, 24, 25, 20, -21, -33, -21, -29, -11, -1, 30, -4, 13, -4, -9, 11, -16, 50, -30, 28, -10, 4, -26, 17, -23, -17, 20, -30, -18, -8, -10, -2, 29, 73, -6, -12, 2, -37, 11, 25, 27, -10, -45, -28, 26, -47, -7, 7, 0, 46, 1, 19, -1, 3, 17, -58, -20, 17, 21, -26, -6, 15, -12, 32, -14, -11, -53, -22, -17, -27, 7, -30, 13, -11, -11, -32, 1, 9, -26, -16, -31, -16, 19, 16, -44, 29, -13, -17, -11, 48, 17, -6, -3, 1, 4, -12, 4, 5, -13, -13, 22, -12, -20, 20, 27, 19, 0, -17, 21, 0, 11, -17, -2, 5, 4, 13, -2, 24, -26, 13, -24, 9, 1, 19, 36, 6, -31, -15, 39, -4, -47, -3, 14, 13, 28, 0, -11, 40, -28, -16, -51, 19, -10, 2, -15, -33, 19, 5, -18, -5, -32, -7, -17, 13, -10, 17, 37, 48, -32, -28, 2, 33, 8, 7, 1, 1, -47, 12, -12, 1, 31, 31, -7, -39, -16, -18, 25, 33, 2, -40, 27, 22, 27, -23, 48, 10, -37, -31, -26, 42, -18, -14, -11, 9, 24, -28, -1, -22, 56, -58, 13, 35, -23, -39, 32, -12, -43, -1, -35, 48, -20, 21, 16, -29, 5, -19, 9, -21, -16, 3, -12, -8, 23, 37, 2, -7, -48, 24, -43, 10, 19, 13, -14, 1, -28, -44, 8, -20, -3, 9, 6, 15, 10, -31, -5, -29, 13, -26, -27, -34, -1, -8, -6, 21, 17, -23, -9, -10, -5, -14, -3, -34, -2, 20, 2, -23, -10, 22, 4, 24, 7, -10, 42, -21, -18, 27, 7, -8, 16, -42, -47, -30, 6, -18, -1, -22, 2, 18, 3, -14, 10, -24, -8, -16, -24, -23, -21, 18, 11, 23, 32, -5, 50, -20, -7, 20, 21, -9, -45, -20, -3, 36, -41, 7, -22, -36, -9, -49, 7, -15, 28, 9, 9, -27, 5, 25, -11, -18, 2, 26, 29, -10, -12, 15, 34, -1, -33, -21, 8, 9, 4, 0, 31, -9, 23, 49, -19, -7, -5, -19, 14, -21, 28),
    (10, 25, 9, 0, -19, -30, -13, 12, 21, 23, 23, -26, 6, -23, 9, 31, 18, -11, -36, -20, -26, 4, 13, -31, 35, -5, 42, 1, -9, -21, -20, 14, -9, -4, 18, -20, -17, 16, 27, -3, -7, -12, 3, -19, -17, -20, 42, 27, 28, -10, 26, -41, -26, 6, 30, 7, 16, -33, 0, 18, 2, 16, 0, -24, -57, -28, 16, -13, -4, 1, -9, -11, -18, 31, -3, 34, 30, 29, 3, -20, 11, -24, 30, -15, -4, -14, -37, 43, 0, -5, -20, 10, 17, -5, 14, -6, -3, 19, 15, 11, 6, -20, -6, 3, -39, 7, -34, 5, -17, 6, 7, -47, 15, -9, 30, -9, -15, -18, -21, 17, 4, 11, 11, -6, -31, 27, -40, -25, 11, -21, 10, 20, -17, -20, 41, 14, -18, 18, -21, 26, -2, 34, 50, -15, -20, 1, -41, 13, -6, 15, -1, 13, 7, 6, 30, -4, -19, -16, 13, -7, -27, -2, -30, -31, -20, -29, -36, 4, -22, -5, 28, -41, -19, 2, 13, 26, -25, -7, -37, 2, -14, 10, 10, -10, 29, 3, -17, 36, 7, -58, -3, 28, -24, -9, -6, 12, 13, 24, 16, 7, 17, 38, -2, 21, 19, -11, 12, -12, -8, 8, -32, 0, -23, -10, 5, -13, 20, -20, -1, -27, -4, 3, -8, -16, 0, -38, 12, 18, -16, -32, -15, 6, 5, 11, -29, 34, 0, -42, -12, 25, 17, -29, 6, -33, 0, 9, 39, 28, -8, -10, -9, 10, 23, 3, -1, 23, -8, 3, 17, -7, 1, 21, -4, -15, 11, -11, 1, 3, 21, 1, 5, -10, -4, -24, -1, 13, 22, 43, -13, 6, 30, -24, -2, -9, 31, -3, -22, -36, -7, 15, -1, 20, -2, -3, 31, -27, -35, -30, -4, -31, -4, -23, 12, 28, 3, -6, -2, -5, 14, -18, -27, -33, -30, -3, -24, 9, 5, -7, 7, -16, -16, 10, -12, -9, 3, 9, -22, -5, 50, 35, 5, 16, -21, -1, 8, -4, 3, 14, -36, -22, -5, 16, 26, -22, 5, 3, 3, 20, -4, -10, 18, -15, -27, 6, 22, 2, 26, 0, 5, -12, 23, -11, 20, -15, 10, -2, -39, 3, 6, 22, -12, 5, 27, 31, 12, -8, -8, -28, 37, 20, 34, 3, -26, 2, 8, -15, -10, 8, -7, 21, 25, -35, 9, -8, 11, -24, 4, 22, 7, 4, 12, -25, 21, 1, -12, -8, 56, 22, 3, 13, 6, -5, -20, 0, 4, -20, -7, 5, 9, 61, -34, 22, 17, 12, 21, -5, 5, -3, -27, 20, -2, 0, -6),
    (-23, 25, -18, 14, 17, 1, -1, -12, -13, -28, 7, 28, -10, 12, -21, 30, -10, -12, 13, 24, -17, 3, 22, 12, -17, 8, 4, -1, 14, 3, 6, 24, -5, 15, -13, -1, -3, 12, -12, -9, 29, -25, 25, -37, -17, -16, 33, -19, -22, 23, -1, 34, -3, 5, -5, -9, 19, 18, -13, -9, -28, 35, 3, -8, 0, -8, 2, -7, -1, -6, 21, 10, 11, 13, -11, 7, -33, -13, -4, 4, -9, 50, 2, 32, 0, -9, -24, -19, 1, -4, -5, 7, 4, -27, 24, -45, 21, 0, -14, 18, 2, 35, -27, 43, 5, 15, 25, -11, -18, 12, 3, -24, -14, -21, 0, -4, -23, -33, 14, -13, 13, 22, -14, 4, -14, 6, 10, 37, -4, 13, -14, 12, 16, -24, -15, -15, 19, -21, 36, -1, -3, -9, 25, -3, -23, -4, -13, 18, 29, -23, 10, 46, -40, -43, -4, 34, -40, -19, 14, -25, -24, 22, 29, -3, -8, -1, 30, 3, 35, 0, 33, -42, -24, 16, 7, 0, -3, 38, -14, -53, 25, -14, 13, -19, 16, -10, -13, -27, -29, -16, -18, 14, 4, 3, 10, 26, -12, -25, 2, 36, 8, -30, -23, 9, -32, -15, 10, 20, -23, -29, 9, -1, -32, 24, 52, -2, 12, 15, 39, -14, -48, 29, 11, 22, -7, 34, -7, -19, 22, -32, 1, -22, -36, 20, 0, -42, 20, -13, 18, 16, -8, -1, -23, 45, 4, -1, -10, 16, -8, -42, 19, 5, -55, -2, 2, 11, -28, -25, 6, -19, 3, 0, 47, -28, 48, -10, -4, 1, -33, 28, -16, 36, -4, 8, 5, 15, 9, -39, 13, -24, -21, -4, -37, -35, -31, -19, 23, 22, -4, 22, -9, 6, 16, -16, -9, 56, 5, -16, -31, -5, -14, -12, -21, -23, 16, 20, 3, 22, 22, 14, -18, -2, 27, 14, 14, -9, -24, 8, 6, 34, 10, 5, -22, -27, 1, -25, -12, 20, 14, 7, -1, -62, 34, 43, -3, -3, 2, 25, -35, 28, 30, -55, -13, 34, -13, 0, -41, 34, 6, -9, -8, -18, -35, -25, 8, -20, -12, -24, -6, -25, 36, 5, 16, 22, -41, -3, -36, 6, 4, -3, 6, -1, 0, -24, 34, -11, -1, -9, -13, -32, 35, -14, -11, -20, -22, 6, -5, 27, 6, -35, 9, 40, -18, -20, 2, 21, -11, -22, 10, -8, 14, -10, -21, -40, -28, -15, 2, -16, 11, -26, -10, 17, -26, -23, 6, 12, -27, -3, -43, -51, -1, -22, -4, 21, 24, 15, -39, -30, -28, -42, -13, 5, 12),
    (6, 42, -9, 4, -8, -26, -43, 2, -16, 10, 14, 31, 16, 4, -27, -46, -20, -11, -19, -6, -20, 20, 32, 15, -7, -11, -27, -14, 26, 23, -16, -13, 6, -11, 19, 10, 11, 40, -3, -16, -44, 19, -5, -3, -23, -9, -3, -8, -12, -23, -17, 16, -2, 31, -23, 10, 6, 25, 15, -12, -23, -29, -12, -26, 0, 27, 1, -15, 37, 20, 18, 20, 13, 43, -16, -13, -12, 18, -1, -19, 21, -15, -7, 28, 24, 7, 3, 8, -16, 10, 2, -4, -32, 14, -25, 24, 25, -20, 9, -2, -34, -10, -15, -18, -5, 40, -22, -1, 15, -25, -12, 3, 21, -6, 17, 7, -7, -28, 21, 32, 29, -1, -23, -21, 19, -17, -22, -5, -4, -34, 2, 9, -15, 7, 31, -23, -25, -27, 5, 13, 13, -23, 4, 12, 0, -14, -16, 7, 19, 10, -36, -19, -17, -24, -49, 16, 7, -8, -23, 5, -11, 9, 14, 4, 18, 1, 18, -32, -11, 24, -24, -52, -11, 28, -9, 28, 6, -25, -14, 17, -24, -26, 34, -28, 33, -1, -13, 10, 24, -33, 9, 3, -1, 8, 6, 4, -17, -17, 17, -12, -21, -22, 12, 48, -12, 18, -14, -36, -26, -38, 16, -30, 3, 31, 44, 2, 40, 35, -32, -36, -28, 36, -6, 26, -24, -32, 35, -8, 2, -4, -4, -28, 5, -42, -17, 25, 7, -14, -43, -7, 10, 22, -18, 0, -37, -13, -28, 38, 29, 32, -34, 22, 9, 9, 2, -5, -1, 18, 11, -25, -8, 26, 33, -1, 31, 21, -26, -2, 6, 22, -46, 18, -31, -2, 16, 15, 23, -4, -1, -11, -20, -30, -9, 0, 15, -8, -5, 7, 9, 23, 28, -20, -15, -4, 2, -4, -10, 3, -19, 17, 31, 20, 2, 14, 16, -16, 2, 22, -18, 8, -21, 1, -29, -16, -44, 3, -19, 11, 8, 8, 16, 0, 27, 6, 11, -15, 0, 0, 24, 15, -28, -3, -16, -18, 18, -15, 15, 20, 31, -3, -14, -39, 22, 22, 22, 13, -3, 10, 7, 11, -19, -31, 1, -18, 5, -5, 13, 1, 11, 25, -4, -23, 3, 38, -27, 25, -6, -24, -14, -31, 31, 27, -30, 19, -14, -26, -11, -6, 6, 4, -31, -35, 1, -23, 8, 57, 18, 29, -20, 9, -31, 40, -25, 10, 0, 2, -18, 9, 6, -3, 4, -23, -32, 3, 16, 1, -2, 12, 11, -26, 13, -18, -1, -12, -28, -9, -27, -3, -24, 16, -22, 25, 4, -37, -9, -2, 13, -3, -6, -12, -15, 18, 2),
    (18, -48, -10, -40, 10, 12, -4, 10, 0, 14, -34, 21, -3, 21, 22, -29, -26, -23, -16, 35, 7, 27, 13, 36, -8, -50, -57, -15, 24, -15, -41, 2, 21, 31, 18, -4, 1, -11, -48, -16, -50, -41, 26, 1, 8, -9, -3, 40, 6, 40, 9, 7, -7, 16, -17, 30, 3, -47, -16, 17, -10, -15, -3, 29, -3, 24, -8, -23, 18, -4, -14, 17, 5, -14, 17, -32, 10, 18, -32, 30, 0, 22, 35, 19, -3, 0, -35, -25, -5, -45, -22, -38, -31, -36, -28, 15, -11, 55, 6, -9, 27, -19, 12, 39, -7, -8, -27, 11, -20, -22, 24, 27, -3, 8, -5, -9, 24, -29, 26, -27, 20, 44, 31, 10, -34, -13, -23, 1, -14, 32, -9, 5, 28, 27, 18, -21, -5, -8, -18, 22, 10, -14, -6, -40, -14, -16, 37, 1, -10, 0, -21, 4, -1, 9, -3, -13, -12, -29, -23, 19, 22, -11, -9, -28, -10, -29, -19, 23, 12, -36, -4, -4, 12, -4, 26, 2, -13, -10, 2, -2, -40, 16, 31, -3, -5, 5, -3, -35, -14, 2, -21, -38, -7, 21, 48, -16, 9, -11, 6, -21, 2, 10, -9, -39, 0, -25, -8, -19, -39, 14, 11, -9, -33, -9, -38, 4, 2, 6, 10, 18, -19, -9, 6, 23, 17, -20, 12, -11, -10, 15, -33, 1, -10, 27, 23, 11, -24, -11, -3, 7, -17, 32, 33, 5, 27, 14, 4, 26, 7, 13, 13, 19, 15, 22, -21, -6, 3, 23, -2, 12, 13, -26, -27, -11, 34, 34, 22, 15, -32, -12, -28, -6, 1, 14, -27, 21, 29, 6, 17, -20, 11, 35, -49, -7, 14, 24, -7, -1, -25, 25, -1, 10, -4, 33, -16, 26, -11, 9, -5, -26, 3, -20, 17, -15, -7, -13, -2, 14, 0, -7, 3, 22, 9, 21, 39, 38, -9, -45, 11, 12, -10, -6, -13, 23, 17, -28, -7, 33, 10, 28, -16, 11, -21, -15, -2, -20, 34, -1, -22, 2, -18, -22, -33, 37, 15, -4, -32, -21, -21, 0, 29, -17, -33, -36, -30, -20, -3, -9, -3, -2, -15, 15, -29, 2, -6, -39, -1, 20, 7, -26, -16, 20, 40, -40, -32, 3, -1, 5, 20, 27, 15, 2, -19, -20, -28, 29, 5, -28, -33, -17, -10, -21, -18, 2, -2, 18, 4, 30, 27, 5, 26, -12, 8, 1, 8, -3, -21, -36, 18, 25, -31, 12, -21, -27, -42, 11, 11, 19, 15, -36, 9, -24, 3, 6, 3, 48, -6, -8, 6, 15, 9, 2, 11),
    (23, -21, -12, 10, -24, 16, -19, 0, 16, -6, -16, -36, -15, -4, -32, 3, 2, -4, 3, -8, -26, -1, 37, 17, -12, -31, -6, -41, 25, -25, 41, -18, -28, -9, 8, -4, -13, -6, -29, -22, 43, 24, 12, -12, -26, -45, -29, 38, 3, -24, -21, -28, 20, -18, -34, -18, -11, -12, 21, -14, -7, 39, -9, -4, 7, -22, -7, 14, 12, -15, 72, 1, -5, -41, -10, -37, 32, -21, 7, -21, -35, -34, -11, 2, -18, 12, 7, -10, 4, 23, 18, -28, 2, 12, 4, 11, 31, -40, -19, 13, 0, -21, -46, -2, -16, -36, 11, -26, -31, 26, -5, -3, 58, 18, -14, 24, 14, 9, 19, 3, -19, -16, -13, -39, 1, -19, 32, -34, 4, 11, 37, 2, 16, -29, 23, -46, -12, 14, 20, 3, -33, -11, 22, 34, -26, -18, 2, -11, -22, -15, -35, -21, -26, -32, -14, -7, 25, 9, -34, -4, 15, -35, 13, 8, 11, 31, 21, 17, -55, 13, -3, -1, 35, 6, 11, 20, 13, 5, 32, -18, -23, -14, -42, 29, 9, 12, 28, -27, -20, -23, -34, 24, -17, -11, -17, -26, -22, 14, -26, -33, -7, -23, -7, -30, 15, 12, -10, -13, 4, -38, -17, 52, 7, 1, 16, 19, -12, -1, -10, 3, -4, -12, 25, -25, -28, -30, 12, 7, -18, 1, -39, 40, 1, 27, 16, -2, -5, -14, 26, 30, -16, -38, -14, 8, -17, 12, -2, -2, 0, -55, 2, 4, 35, -6, -37, -7, 7, 21, -27, -13, -18, 12, -5, 34, -56, -25, -9, -1, -8, -31, -41, -19, -42, -12, -4, 19, -6, 3, 8, 25, 45, 5, -4, 13, 7, 12, 48, -1, 3, 26, 12, -12, 29, -15, -9, 1, -25, -5, -13, 8, 0, -12, -7, -4, 20, -25, 27, 3, -12, -7, 19, -20, 14, 12, 18, -6, -23, 22, 23, -12, 16, -53, 26, 27, -39, 17, -9, 26, 30, 12, 33, -17, -7, 3, 2, 14, 0, -18, -29, -17, 19, 13, -4, -26, -9, -15, 1, -3, 31, -1, 32, 8, 42, -9, 19, 38, 32, 21, 6, 18, 10, 18, 6, -17, -6, 2, -46, -23, 3, -35, -2, -6, -35, 13, 9, 15, -2, -35, 24, -15, 8, 37, -21, 19, -4, -8, 33, -10, -7, 18, -26, -42, -19, -5, 18, 5, 0, 0, -26, -13, 64, 17, -6, 13, 33, -37, -19, -2, -8, -23, -10, 28, 22, 11, -16, -18, -35, -5, -9, 32, -47, -2, 48, 8, 8, 5, 9, -12, -1, -4, 50, -24, 16),
    (17, -41, 4, 40, -6, -5, -15, 36, 30, -11, -11, -14, -20, 2, 14, -51, 46, -14, 27, -36, -30, -19, 24, 29, 20, -35, -52, 15, 4, 13, -40, -16, -66, -29, 21, 17, -8, 12, 12, -17, -5, -35, -32, 6, -39, 8, -11, 10, -13, -50, 18, 33, -11, -9, -3, 15, 30, -21, -24, 8, -7, 4, 4, -32, 5, 13, -17, 12, -6, 6, -11, -7, -4, -33, -18, -21, -11, 22, -16, -32, -47, -14, -19, -25, -17, 51, 4, -6, -21, -20, -26, 15, -22, 29, -4, 21, 13, -33, -16, 53, 17, -1, -8, 1, 0, 23, -7, 40, -32, 4, 26, -8, -18, 15, 0, -1, -1, -3, -9, -22, -1, -2, -22, -29, 11, -11, -35, -47, -28, -8, -12, -12, -27, 10, 41, 7, -29, -37, 2, 55, 13, -3, -13, 20, 10, 44, 9, 13, 6, -18, 27, 13, 0, 46, -50, -24, 39, 17, -35, 14, -24, -1, 16, -8, -45, -36, -3, 17, -18, -31, 22, 30, 31, -10, -42, -28, -1, -21, -32, -34, -20, 3, 10, 11, 13, -6, 14, -20, -19, 21, -10, -16, -23, 18, 12, -28, 10, -24, 22, 42, -24, 18, -14, -37, -12, 33, 16, 6, -10, 13, -9, 17, -25, -49, -31, -8, -17, -42, 24, 35, 18, -6, 9, 17, -8, 17, -3, -8, 11, 1, 12, -4, 7, 9, 4, 26, 18, 20, -12, -36, 3, 16, 15, 12, 28, -9, 22, -6, 25, 24, 2, -12, 18, 13, 12, -11, -37, -28, -6, 24, -8, -26, -13, 0, 29, -28, 8, 27, 19, 8, 15, -26, 3, -13, -14, 21, 29, 19, -4, 16, -12, 35, -23, -8, -38, -8, 0, -14, 0, 1, -5, 13, 8, -20, 9, 5, 4, -5, -8, -26, 14, 31, 19, -34, 3, 16, -19, 8, 3, -4, -9, 6, -19, 13, -14, 17, -36, -34, -16, -5, -3, 2, -22, 14, -10, -8, 15, 11, 33, -16, 19, 21, -6, 28, 2, -21, 2, -28, 24, -31, 20, -30, 20, -16, 22, 3, -11, 6, -9, 24, -11, -21, 25, 4, 12, 6, 16, -18, -61, -1, -24, 0, 7, 1, -17, 4, -48, 15, -8, -9, 14, -8, -8, -6, 8, 34, 17, 14, -9, 46, -14, 26, -21, -28, -28, -10, -23, -4, 10, 13, 5, -14, 17, 15, 21, 8, -13, 11, 5, -17, -26, 5, -21, -10, 11, -8, 8, -34, 19, 2, -5, -20, -30, -5, 4, -6, -1, -26, 8, -34, 27, 15, 13, 31, 34, 33, -11, -3, -26, 29, 30, 21, -13),
    (-13, 16, 17, 3, 24, -21, 18, 21, -26, -20, -29, 26, 15, -24, 11, 1, 6, -44, 12, -16, -14, -4, -29, 2, 37, -21, -15, 24, -13, 14, -14, 15, -4, -7, 0, 7, 10, 25, -16, 7, 5, 7, -36, -26, -32, 12, -25, 18, -29, -4, 45, 3, 4, 13, -4, 14, -31, -23, -31, 26, -51, -31, 27, 19, 9, 8, -17, 12, -2, 26, 14, -31, -10, 18, -9, -8, 3, 13, 2, -35, 23, 8, -25, 10, 16, -9, 6, 13, 15, -24, 9, -35, -6, 0, 6, 7, -13, -22, -21, 0, -11, -12, 8, -26, 30, -24, 4, -35, -10, -12, -15, -6, 2, 8, -34, 28, 13, -22, 48, -29, -12, -15, 47, 8, -30, -23, 21, -10, -33, 16, 12, 8, -12, 2, 40, -13, 6, 19, 3, -21, 0, -6, -21, 22, -12, -3, 20, -11, 6, 9, -2, 34, 22, 41, 12, 3, -1, -24, 1, -2, 49, -4, -17, 21, 8, -19, -30, 22, 23, -3, 24, 31, 9, -28, -17, 25, -7, 20, -11, -5, 19, 22, -21, 27, 12, -2, 29, -22, 17, -27, -12, -21, -29, -8, 54, -34, 12, 6, 48, 23, -12, 33, -4, -5, -2, -15, 29, 45, 32, -5, -28, 11, -47, -3, -8, -27, 32, 6, 11, -9, -12, -6, -1, -24, -24, 20, -28, -1, -16, 37, -4, 12, 3, -26, 50, -2, 32, 1, -1, -22, 15, -3, 42, -4, -19, 1, 4, 15, 12, 33, -8, -5, -5, -33, -16, 23, 18, 4, -25, 3, -29, 5, -5, 18, 3, -22, 26, -13, 41, 4, -13, 4, -16, 24, -19, 19, 12, 12, -1, -14, -20, -10, 41, 7, 1, 7, -12, -4, -17, 12, -30, -23, 7, -14, -1, -25, -18, 11, -18, -30, 54, 7, 9, 5, -20, -4, 5, 5, 8, -27, -15, -6, -34, -18, -11, 35, -17, -44, 6, 2, -7, -24, 3, 10, -19, -13, 11, -2, -7, 27, 4, -27, 4, 10, 21, -11, 14, 5, -27, 17, -21, -12, 21, 6, 3, -1, -23, -13, 12, 7, 31, -20, -24, 0, 12, 21, -1, 5, -31, 19, 29, 48, -22, 4, -4, -26, -3, 3, -6, 6, -26, -20, -23, -17, -16, 25, 9, 10, -24, 17, 25, 7, -32, -19, 17, -7, -61, -13, -29, -5, 7, -26, 6, -2, -3, -32, 1, 5, -4, -18, -29, -27, -15, 21, 0, 5, -10, -8, -18, 35, 11, 19, -17, -15, -3, 7, 7, 18, -14, -42, 14, 20, -32, -11, 34, -5, -24, -28, -24, -15, 15, 18, -10),
    (23, -15, 23, 10, -16, 10, 4, -51, -3, -6, -7, -6, -53, 0, 12, -29, -34, 24, 2, -14, -26, -23, 1, 8, -6, -15, 23, 6, 13, 21, 15, 20, -7, -12, -2, -1, 43, 31, 1, -42, 21, 18, -12, -9, -26, -20, -12, -24, -36, -16, -18, -34, 29, 7, -23, 14, 8, -7, 30, -4, -3, 0, -7, -13, 16, -6, -28, -16, -11, -2, 27, -1, -3, 19, 7, 0, -25, -22, -15, 0, 16, 26, 13, -7, -29, -17, 24, 8, 2, -31, -8, -19, 8, -10, 20, 8, -9, -59, -28, -7, -5, -26, 6, 9, -22, 2, 20, 13, -34, 13, -7, -20, 43, -5, -4, -6, -16, 34, -3, -8, 2, 32, 16, 8, -35, -19, 4, 17, 9, 16, 31, -26, 9, -23, 12, -37, 2, 6, 36, 28, -24, 4, 12, 32, -2, -11, -21, 34, -23, 6, 5, 17, 26, 17, -6, -36, -42, -28, 18, 8, -14, 1, -38, -10, -15, 3, -8, -53, 10, 4, 5, -28, 15, 3, -7, -23, -27, -17, -12, 18, 10, -35, 15, 20, 25, 25, 27, 26, -14, 19, -30, -32, 0, 16, 16, -3, -37, 11, -21, 7, 34, 43, 30, -18, 9, 2, 22, 24, 5, 23, -40, -6, 2, 7, -16, -37, -23, 26, -1, 4, 18, -16, 20, 11, -2, -22, -8, -4, 9, -27, 22, 29, -8, 9, 8, 4, 3, 26, -4, -6, 18, -41, 29, 17, -37, -9, 16, -13, -6, 39, 11, -6, -29, -9, -23, -6, -5, -31, 6, 11, -12, -3, -19, 0, -6, 5, -15, 4, -22, 36, 18, -12, -10, -36, -20, 14, 7, -26, -25, -26, 7, 12, -6, 3, 20, 16, 23, 18, -48, -33, -10, 2, -3, 2, 14, 2, 28, 20, 19, -17, -14, -18, -44, 8, 3, -7, 19, -26, -12, -10, 36, -29, 1, 14, -19, -3, -4, -12, -24, 12, -33, 17, 3, -28, -34, 24, 11, -3, 39, 8, 31, -19, 27, -38, 13, 8, -37, 26, 14, 2, -17, -12, 24, 21, 3, -7, 34, -7, -19, -33, -9, 11, 27, -2, -20, -22, 0, 6, 34, 11, 5, -10, 44, -6, 12, -10, -58, 8, -15, 14, -22, 21, 13, -9, 9, 0, 16, 35, 29, 22, -13, -1, 47, -13, -32, 10, 15, -16, 1, 24, -12, 43, 13, 17, 30, 1, 17, 1, 12, 23, -12, 20, -41, -30, 10, 13, -27, -28, -15, -9, 7, 2, 31, 17, 18, -17, 16, 13, -16, 37, -19, 8, -17, 6, -8, 11, 9, -10, 17, -36, -16, -26, -4),
    (-39, 28, 23, -36, -7, 31, -22, 11, 15, -1, -42, 19, 19, -5, 10, -17, -13, 16, 11, -32, -16, 21, -21, -1, -13, -15, -38, 6, -8, 22, -27, 26, 21, -12, -13, 9, -29, -42, 0, -31, -5, 20, -24, -7, 4, -14, -6, -33, -30, 53, 10, -12, 16, -11, -24, 34, 2, -2, -10, 33, -19, -13, -2, 14, -31, 2, 27, 4, -18, 20, -11, 11, 46, 2, -2, -37, -11, -2, -8, 27, 33, 22, -13, -1, 29, -36, -11, 15, 2, 23, -11, 15, -19, -3, 7, -23, -16, 28, -22, 15, 14, 15, -9, 20, 14, 4, -13, -8, -24, -28, 24, 8, 5, -8, -4, -8, -4, -8, -28, -17, -30, -2, -24, 6, -52, 4, 24, -13, -16, 42, -36, -31, -10, -65, 14, 14, -26, -7, -37, -21, -9, 3, -29, 14, 2, -13, -2, 6, -31, -5, 0, 10, 4, 11, -12, -13, 16, 36, 21, 13, 13, -13, 3, 21, 22, 31, -19, -30, 14, 15, -14, -5, -18, -41, -45, 6, -18, -15, -23, -18, -15, -17, -30, -8, -7, 12, 9, -8, 0, 9, -8, -5, -15, 16, -12, -55, -10, -33, -2, 33, -25, -27, -25, 1, 5, 10, 6, 5, -34, -17, -9, -24, -27, -14, 32, -27, 20, 8, 11, -22, -31, -23, -6, 31, -11, -24, 22, 7, -6, 14, -6, -10, -9, 5, -33, 10, 18, 35, 22, -38, 11, 27, 11, 29, 1, -34, -4, 44, 12, 25, -29, 21, -4, -14, 10, 0, -11, 25, -12, -10, -23, -18, -27, -26, 20, 34, -24, -6, 4, -9, -46, -11, -15, -15, 4, -25, 12, -18, 19, 25, -21, -21, 6, -6, -3, 19, 19, -9, -27, -10, 17, -27, 0, 2, 10, -19, 2, 29, 29, -25, 35, -14, -4, -19, 6, -15, -2, 16, -9, -12, -1, 13, -20, 8, -25, -29, -13, -2, 19, 10, -21, -28, -10, 27, -60, 24, -11, -26, -10, 7, 39, 50, -5, 43, 9, -3, 32, 12, 12, -27, -5, 23, 12, -25, 5, -21, 21, 4, 25, 9, -10, -11, -13, 6, -1, 46, -10, 3, -30, 9, 14, -3, -23, -18, -4, 16, -19, 24, 6, -7, 5, 50, 10, 9, -13, -14, 2, -26, 23, 13, -5, 7, 6, 24, 1, 13, 14, 23, -29, 25, -17, 31, -19, 26, -14, -27, -17, -6, 31, -14, 35, -21, 17, 20, -11, 12, -2, -1, 17, -25, 12, 25, -16, 17, -7, -1, -12, -26, 17, 21, -29, -7, 55, -14, -16, 17, 9, 13, -9, -6, 4, 21, 6),
    (2, 5, -7, 17, 22, -9, -5, 23, -33, -4, -37, 37, 15, -15, 15, 5, -7, 4, -5, -24, -21, 13, 25, -7, 44, 0, 30, -13, -20, 35, -1, 11, -19, -6, 16, -33, 15, 45, 0, 4, -15, -3, 10, -8, 33, -4, -26, -43, -16, 41, 13, 24, 2, 29, 5, 6, -16, 24, -29, 0, 3, 14, -25, 18, 30, 31, -19, -29, -24, 31, -1, -6, 10, -23, 19, -18, -17, 19, -5, -8, 28, -9, -19, 29, -15, 1, 0, 1, -12, 29, 20, -1, 34, -6, -39, -51, 8, 24, -8, 13, 6, 4, -19, -3, -28, 33, -30, 13, 22, -7, 32, 14, -4, -17, 10, -45, -10, 22, -34, 32, -5, 26, 9, 19, -13, 1, -25, -13, -14, -11, -11, -19, -6, -2, 37, -10, -28, 30, 6, -22, -19, 4, -17, -57, 27, -16, 0, -50, -15, -13, 12, -9, -10, -29, 10, 25, -17, -16, -6, -17, -29, -7, -31, 2, 2, 12, 59, 5, -26, 0, 17, -18, 22, 11, -18, -13, -32, -12, 35, -3, 22, 61, 0, 8, -25, -17, 45, 14, 40, -10, -12, 2, 13, 5, -2, -29, 4, -19, 3, -5, -24, -40, -2, 16, -29, -35, -6, -35, 8, 32, -27, -34, 26, 22, 28, 10, 30, 27, 2, -28, 21, 13, 0, 21, 17, -10, 32, -31, 32, 12, -24, -8, -44, -24, 25, -24, 4, -29, 6, -22, 21, 3, -22, 1, -7, -27, 13, 16, -9, -40, -8, -9, -40, 13, 35, -24, 32, 16, 31, -22, 8, -19, -3, 23, 4, 6, -19, -34, -8, -8, -25, 4, -14, -19, -2, 1, -33, 9, 16, 1, 0, -52, 19, -29, 1, -33, -7, -2, 13, 3, 6, -1, -13, -6, -27, 12, -1, 12, 20, 27, -8, -8, -34, 26, 8, 7, -11, -6, -9, 13, 55, 7, -19, -9, 28, -8, 8, 17, -5, 1, -20, -20, -19, 16, 1, 11, 17, 0, -39, -7, 6, -2, 31, -29, 0, 26, 40, 1, -13, 4, 17, 3, -21, 15, -27, 15, -7, 18, -2, 8, -16, -29, -33, 31, 18, -27, 25, -11, 12, -22, -6, 7, 13, -12, 1, 0, -3, 11, -31, -20, 5, -40, 21, 6, 18, 26, -7, 9, 6, -29, 2, 14, 33, -11, -12, 9, 8, -23, 11, -13, 25, 16, 10, -12, 18, 8, 31, -1, -10, -4, 25, -17, 5, -1, -19, 16, 21, 4, 41, 4, -23, -8, 0, 11, -11, -1, -18, 11, -13, -54, -3, 12, -5, 11, 14, -5, 7, -3, -8, -11, -13, 14, -1),
    (-1, 9, 21, -63, 6, -38, 5, 17, 11, -25, -27, 38, -9, 13, -26, 3, -8, 2, 29, 13, -11, 3, -51, 22, 5, -22, -12, 17, -19, 0, 18, -5, -7, -13, -12, -22, -37, 40, 3, -5, -24, -1, 1, -31, -13, -43, -17, 13, -28, 0, 18, 51, 0, -8, -30, 21, -18, 23, 7, -8, -22, -34, 3, 12, 59, 11, 21, -4, -72, 11, 38, -10, 39, -11, -11, 21, -46, -1, -1, -5, -10, 30, -21, 31, -9, 2, 29, 3, -11, -9, 5, 15, -10, 9, 7, -6, -4, 44, 35, 10, -13, -9, 19, 21, -22, -9, -27, -18, 21, 28, -4, 18, 21, -11, 13, 24, -45, -4, -16, -23, -27, -21, -20, 27, -22, -33, 22, 10, 14, 11, -2, 31, -17, -9, 9, -27, -18, -27, 0, -20, -4, -24, -7, -7, 5, 26, 26, -7, -10, 30, 9, -16, -10, -18, -7, -28, -41, -23, -43, -20, 9, 46, -27, 6, -9, -8, -15, 14, -3, 6, 44, 0, -37, -11, -1, 30, -17, -20, 35, -3, 4, -3, -13, 45, -33, 31, 12, -41, -7, -40, 3, -38, -26, 32, 40, 27, 18, 17, 0, 16, 1, 15, -16, 13, -14, -35, 3, 10, 31, 8, -24, 4, -8, -36, -2, 7, 34, 11, 37, 45, 0, 13, -6, 13, 5, -22, -33, 23, 13, 32, 43, 27, -8, -12, -6, -22, -5, 14, 8, 0, 7, 7, 40, 0, -19, -21, 28, 29, -11, 49, 17, 9, 1, 20, 39, 44, -1, -48, 0, 32, -3, -11, -23, 1, -4, -33, 23, 10, -18, 50, -25, -10, 13, 27, 12, -20, 11, 8, -13, -31, 10, 11, -20, -17, -7, 20, 1, 4, -8, 36, 14, 9, 5, 36, -8, 0, 37, 23, 1, -8, -23, -4, -7, 36, -10, -9, -4, -7, -11, 16, 6, -29, -1, 14, -7, 9, 21, 24, -27, 0, -10, -4, 38, 21, 7, 7, 24, 23, -16, 3, 25, 28, -11, -8, 8, -32, -31, 23, 12, -8, 17, 1, -33, 16, 30, -9, -22, -23, -8, -12, 26, 34, -6, -2, -16, 2, -23, 27, 15, -7, -31, -7, 1, 26, 5, 22, -44, -12, 1, 21, 0, -29, -4, 1, -11, 20, -21, 15, 19, 22, -6, -13, 11, -31, -7, -7, 10, -39, -10, -1, -22, -6, 2, 14, -15, 18, -7, -7, 4, 21, 19, -24, 15, -6, 19, 15, -5, -11, -2, -33, 11, -14, -13, 13, 9, 44, 1, 25, 21, 21, 34, 0, -18, -19, -8, 12, 24, -27, 5, -30, -11, -5, 11),
    (0, 2, -11, -48, 14, -2, -17, -35, 3, -21, 14, 6, 7, -10, 15, -7, 10, 21, -18, 5, -4, 15, 12, 29, -33, -38, -6, -15, -11, -12, -2, 3, 16, 16, 13, 22, -12, -1, -4, -5, -3, 1, -13, -12, 14, -30, 26, 39, 4, -12, 7, 21, -18, -3, -23, 12, 22, 15, 3, -22, 28, 7, -4, 18, 62, 37, 18, -10, -15, -35, 12, -7, 0, -16, 1, 18, -32, 25, 25, 29, 17, 14, -24, 18, -23, -15, 15, 27, -34, -8, 42, -40, -24, 1, -2, 19, -47, 39, 10, 24, -11, 9, -23, 31, 4, -29, -37, 7, 30, -3, -33, -5, 3, 28, -3, -12, -47, -34, -4, 27, 25, -37, 14, -1, 27, -13, 24, 14, 18, 40, -14, 17, -10, 5, 9, -12, -7, 2, 43, -28, -7, -15, 10, 31, 3, -1, -9, 12, -4, -37, -14, -13, 8, -17, -29, -7, -20, 14, 26, 3, 21, 30, -30, -8, 10, -22, 31, 6, -2, 0, -9, 5, 0, -17, 30, -19, 24, 36, 5, 11, 9, 13, 21, -37, 0, -35, 1, -26, -35, -9, 32, 59, -18, -16, 4, 48, -12, 0, -26, 41, -19, -32, -4, -5, 7, 1, -28, 5, 24, 28, 10, 22, -14, -3, 33, 6, 51, 4, 2, 39, -18, -40, 31, -23, 2, -2, -16, 7, -21, -3, 20, -23, -1, 8, -47, -45, -9, -7, -2, -9, 4, 8, 1, 1, 9, -11, -7, 21, -31, -14, -24, 9, -1, 10, 36, -30, 15, 31, -14, 5, -11, -53, 4, -30, 16, 10, 6, 17, -7, -11, 0, 14, 22, 7, -60, -3, -10, -47, 26, -23, 11, -4, -8, 4, -32, -24, 30, -19, -13, 22, 12, 30, 9, -45, -27, 10, -22, -25, 24, 10, -47, -23, 12, -18, 15, 52, -9, -45, -14, -28, 18, 7, 15, 5, 34, 35, -6, -12, 7, 0, -18, 23, -27, -7, 5, -1, 11, -28, 25, 7, 1, -21, -22, -25, 10, 27, 43, -5, -4, 13, -30, -6, -25, 25, 35, -14, 26, -12, -11, 6, 16, -28, 17, 45, -6, -16, -31, -49, -1, -25, 15, 18, 12, 10, 23, 0, 9, -17, 14, -17, -38, -14, -21, -1, 22, -1, -24, 36, 39, 7, -25, -35, 1, 16, 14, -7, -23, 1, 8, 14, 18, -1, 15, -8, 22, -27, 3, 19, 21, -10, -39, -5, -7, 0, -5, 8, 11, -17, 25, -5, 12, -14, -15, -6, -16, 16, -18, -35, -30, -3, -1, 4, 9, -16, 17, -18, 2, 9, 25, 14, -10, 21, 9),
    (-34, 32, -22, -22, 19, 11, 1, 13, -2, 16, -8, 11, -17, -23, 18, -6, -23, 38, -1, -10, -10, -14, -47, 21, 28, -17, 17, 15, 12, -40, 2, 9, -16, 27, 6, -8, 34, -5, -4, -9, -14, 5, -37, 2, 8, 7, -12, 15, -12, 30, 5, -32, -1, -38, 27, 1, 5, -38, 28, 6, -48, -23, -2, -14, -17, -19, -8, 1, 27, -19, -12, 10, 29, -9, 26, 0, -40, 0, -24, -9, 10, -18, 34, -30, 16, 30, 8, 8, 27, -9, -12, -21, 8, -25, -11, 25, 13, 0, -23, -2, -12, -26, 27, 9, 34, 8, -12, 11, 8, -10, 10, 25, -7, 14, 7, 15, -16, -28, -28, -31, 26, 22, 38, 35, 22, 6, 10, -5, -5, 15, 39, -27, 3, 9, 15, 10, 14, -7, 12, -10, 4, 4, -1, -17, -22, 19, 17, 15, -14, 4, -26, 7, -30, 3, 20, -16, 15, -1, 16, 24, 33, -28, 7, -23, -22, -24, -6, -33, 33, 9, 11, 39, -16, 9, -28, -17, -33, 44, -24, -6, -2, -5, -24, -20, -7, -19, 7, -20, 9, -10, -27, 19, 35, -6, 0, -27, -11, 29, -2, 12, 12, -36, 9, 2, 1, 15, -2, 7, 34, -11, 12, 9, 10, -14, 31, -16, 25, 14, 22, 10, -14, -15, -47, 31, 11, -8, 36, 4, 29, 9, -11, 9, 9, -42, 15, -22, 14, -22, -3, -11, -13, -22, -32, -20, -5, 15, 20, -32, 19, -27, 6, -5, -35, 1, 8, -24, -6, -19, -20, 5, 16, 4, 22, 20, 20, 18, -6, 4, 21, -3, -46, -1, -27, -28, 30, 8, -12, 5, 8, 9, 6, -19, -27, -13, 22, 20, 30, 30, 36, 10, -42, 43, -2, -29, 29, -4, -5, 14, 11, -5, 34, -2, -17, -16, -16, 4, -33, -6, 31, -27, -1, 2, 33, 21, -7, -28, -27, -32, 5, -38, -15, 2, -3, 1, -6, 38, -47, -17, -17, -30, 3, 6, 40, 26, -44, 3, 32, -6, 1, -1, -5, 13, 5, 20, -1, 2, 8, 29, -25, 0, -18, -22, 13, 40, -29, -10, 31, 10, 13, 15, 36, 5, 0, 27, -9, 14, -4, 8, 0, 10, 8, 7, 18, 17, 20, -11, 18, -28, -2, -26, -3, -30, -38, 21, -2, -17, 23, -12, -34, 7, -7, 3, 30, 41, -27, -28, 10, -12, -2, -1, 17, -23, -32, -17, -7, -27, -4, -31, -18, -8, -11, 24, -24, -3, 10, -17, 10, 12, 0, -12, 10, -1, 21, 11, -19, -7, -14, 8, -3, 11, -9, 5, -12)
  );
  ----------------
  CONSTANT Flatten_1_Columns : NATURAL := 4;
  CONSTANT Flatten_1_Rows    : NATURAL := 4;
  CONSTANT Flatten_1_Values  : NATURAL := 48;
  ----------------
  CONSTANT NN_Layer_1_Activation : Activation_T := relu;
  CONSTANT NN_Layer_1_Inputs     : NATURAL := 768;
  CONSTANT NN_Layer_1_Outputs    : NATURAL := 10;
  CONSTANT NN_Layer_1_Out_Offset : INTEGER := 4;
  CONSTANT NN_Layer_1_Offset     : INTEGER := 0;
  CONSTANT NN_Layer_1 : CNN_Weights_T(0 to NN_Layer_1_Outputs-1, 0 to NN_Layer_1_Inputs) :=
  (
    (30, 8, 3, 5, -9, 7, -22, 5, 8, 6, 9, 6, 8, -13, -4, -2, 11, -17, 6, -26, -37, 1, 1, 0, -13, 22, -4, 4, -12, 2, -9, -17, -34, 11, 8, -6, 32, -1, 9, 9, -12, -9, -9, 6, 18, -12, 2, 9, 24, 2, -7, 5, 11, -15, -4, -2, 23, -15, 6, 8, 0, -4, -16, -5, -1, -2, -13, -12, -24, 16, -3, 10, 22, 29, -2, -16, -22, 6, -3, -2, -22, -1, 0, -8, 20, -2, 13, -1, 18, -9, -23, -17, 7, -24, 9, -19, -8, -11, 2, -3, 22, 2, -31, -17, 16, -16, -3, 13, 9, 6, -12, 10, -6, -2, -17, -2, -31, 23, -2, -11, 6, 10, -7, -11, -1, -2, -23, 7, -18, -2, -5, 8, 12, 7, -1, 5, -2, -4, 2, 0, -13, -23, 21, 11, 2, -3, -3, -6, 10, -16, -14, 13, 14, 2, 7, 9, -12, 5, -2, -13, 5, -1, -3, 3, -12, 5, -14, -14, 18, 12, -13, 1, -11, 2, -35, -4, -7, -6, 9, -1, 21, 10, 1, 4, -5, -16, 15, -2, -4, 0, -7, 4, 15, -18, -2, 9, -5, 1, -46, 6, 7, 10, 28, 11, 14, -17, -9, 12, 12, -8, 0, -20, -20, 27, 20, 13, -7, 15, -8, -7, -5, 7, -13, -6, -24, 14, 21, -19, 18, 0, 6, 13, -2, -28, 0, 6, -11, 22, 15, -8, -17, -16, 5, 4, 6, -12, -13, -14, 26, 0, -1, 8, -9, -18, -17, 9, -32, -47, -9, -20, -47, 15, 14, 6, 0, 12, 10, -15, -12, 19, -10, -29, 4, 9, 2, -8, 3, 0, 10, 14, -4, -16, -15, -14, -14, 19, 13, -11, -3, -16, 9, -8, 21, -3, -12, 2, 22, 11, -23, 12, -2, -11, -24, 11, -24, -13, 9, -18, -50, 8, -14, 11, -7, 1, 18, 10, -18, 25, -19, -19, 1, 3, 8, -11, 10, 14, -6, 5, 3, 6, -20, -1, -34, 1, 1, 7, -7, -18, 6, 5, 13, 0, 3, 5, 27, 7, 2, 16, 7, 0, -20, 14, -11, -2, 7, 7, -30, 10, -16, -10, 9, 17, 4, 22, -12, 3, -1, -10, -18, 11, -9, -5, 17, -5, 6, 4, 20, -18, -9, -5, -2, 1, 0, -13, -9, -10, -3, 5, -8, 10, -23, -18, 22, 6, 18, 10, 9, -18, -5, 14, -1, -35, -10, -20, -5, 26, 18, 6, -17, 21, 2, -10, 8, 29, -30, -9, -32, -8, 21, -26, 3, -22, -13, 14, -36, -34, -2, 18, -5, 32, 15, -19, 0, -29, 6, -22, 15, 0, -7, -16, 17, -6, 13, 11, 1, 2, -4, 12, -24, -46, 8, -15, -4, 15, 18, 3, -11, 21, 3, 7, -1, 17, -22, -20, -10, -6, -4, -10, 2, -7, -3, 11, -4, 1, -19, 0, -7, 8, 20, -14, -12, -21, 14, -16, 14, 9, -8, -1, 15, 12, -1, 4, 11, 6, -15, 13, -27, -22, 5, -19, -8, 3, -5, 14, -6, 19, -11, 3, -18, 37, -6, -17, 2, 9, 14, -22, 5, 1, -4, 24, 1, 8, -9, -7, -12, 29, 13, -5, 1, -1, 7, 9, -1, -15, 10, 0, 10, 19, 5, 9, 4, -6, -10, 3, -15, 0, 4, -6, 0, -4, -21, -6, -2, -6, -21, 16, -5, 0, 0, -14, -1, 2, 3, 11, 5, 19, -4, 9, -3, -3, -4, -1, 1, -8, -1, -5, 3, -22, -2, -20, -4, -6, -10, -7, 28, 6, 16, 1, -2, -12, 5, 10, -3, -45, 2, -22, 3, 8, 11, -17, 1, 13, -3, 12, 7, 4, -23, -4, -21, 4, 3, -8, 5, -16, -26, 8, -20, -1, -1, 3, 6, 17, 9, -6, 3, -29, 9, -16, 13, 2, -7, -13, 2, -7, 13, 1, -7, -10, 6, 7, -10, -43, 7, -13, -12, 8, 4, -11, 7, 28, -10, -1, -5, 9, -22, -15, -1, -1, 11, -4, 4, -2, -24, -7, -6, -15, -9, 1, -5, 18, 6, -4, -3, -27, -1, -3, 12, 0, -11, 18, 16, -6, 0, 3, -1, -9, 7, -8, -29, -11, -2, -1, -5, 8, 2, 1, -3, -1, 2, 0, -12, 26, -6, -7, -2, 26, 5, 11, 4, 8, -14, 6, -2, -11, -7, 12, -8, 4, -1, -17, -6, -6, 9, -3, -1, -5, 2, -3, 21, 2, 6, 8, 1, -16, 12, -8, -12, 0, 8, -20, -13, 10, 3, -5, -4, -5, -18, 7, -2, -4, -4, -16, 13, 19, -9, 10, -12, 3, 6, 0, -10, -5, -1, 1, 5, 23, -10, 8, 5),
    (22, 14, 10, -9, 8, -22, 0, -7, 14, -6, 16, -32, -17, -17, -19, 11, 5, 20, 19, 22, -5, 3, -7, 10, -20, -14, -7, -4, -20, -19, -6, -6, -4, 9, -16, 4, -9, 16, -6, -5, 5, -4, -22, 13, -1, -12, -1, 10, 1, 12, -15, 9, 13, -7, 9, -18, 5, -15, 11, -48, 15, -1, 1, -19, -7, 12, 35, 3, -16, 13, 14, 9, -20, -5, 8, 6, -18, 3, -6, -16, 1, 2, -3, 7, -21, 12, -29, 9, 13, 17, -33, 3, -18, -21, 5, 4, 8, -12, -9, -4, 14, 12, 5, -8, 5, -17, -13, -20, 6, 4, -1, 6, -23, 9, 40, 13, 5, 13, 10, 4, 8, -7, 2, 5, -7, -9, -5, -6, 12, -9, -2, -11, -27, 6, -9, -1, -9, 23, -26, 17, -14, -22, -22, -9, -2, -19, -5, 9, -4, -2, -11, 11, 7, 0, -17, -14, -8, 7, -3, 8, -3, 5, 12, 14, 5, -6, -3, 17, 10, -5, 0, 9, -26, -2, 1, -3, -4, -5, -4, -14, -6, -1, 12, -8, -3, -3, -15, 10, 8, -14, -9, -20, -19, 15, -1, 18, 7, 13, -9, 1, -5, -1, -23, -24, -4, -1, -5, -11, 4, 23, 11, 10, 3, -9, 5, 0, -9, -33, 13, 21, 14, -9, -27, 6, -8, 18, -20, 13, -20, 5, -9, -17, 13, -15, -23, 1, -20, -14, -14, 5, 7, 6, 12, 12, 19, 17, -2, -23, 0, -5, -7, -21, 14, -8, 8, 1, -13, 4, 16, 9, -4, 16, 17, 17, -12, -32, 13, 0, 15, 15, -13, 3, 15, -1, -26, 8, -20, 12, 22, -2, 8, 6, -24, -10, -23, -5, -2, -6, 8, -7, 13, 25, 15, 12, -5, -11, -2, -17, -18, -11, 6, -16, 9, -11, -20, 15, 21, 5, -11, -5, 1, 14, -13, -42, 14, 14, 4, 3, -7, -12, 19, 5, -34, -13, -33, 5, 27, -6, 13, 7, -11, 0, -16, -4, -5, 8, -6, -2, -12, 29, -2, 3, 2, -4, 15, -4, -6, -17, -1, -18, -6, -2, -24, 4, 11, 14, -24, -29, 2, 13, -2, -19, 6, 4, -9, 2, -7, 0, 9, -5, -21, 0, -23, -16, 33, -5, 28, -2, -24, 6, -2, -10, 3, -4, 12, 21, -19, 2, 8, 12, -7, -16, 4, 16, -15, 4, -4, -11, -5, -8, -12, 12, 1, -9, -7, -11, -1, 2, -7, -5, 0, 6, 9, 4, -15, 17, 3, 9, -10, 1, -2, 9, -1, -6, 2, -11, 1, -28, -14, -6, 2, 12, -7, -5, 3, 18, 6, 5, 11, -12, 6, 4, -4, -4, 0, -10, 7, -3, -5, 12, 13, -1, -10, -13, 13, 1, -8, -14, 5, 12, 3, 11, 5, 10, 11, 1, -24, 11, -16, -2, 0, -15, 9, 9, -10, -24, -16, 1, 13, 8, 11, 2, -4, 18, 1, -6, -2, -15, 10, 6, -7, -9, -2, -9, 7, -4, 3, 10, 10, 9, -3, 0, 0, 8, -5, -26, 6, 8, 8, 1, -1, 10, 16, 26, -34, 14, -18, -2, 19, -8, 19, 3, -21, -22, -5, 2, 9, -6, -7, 1, -12, 13, -2, -1, -5, -10, -4, -7, -14, -10, -9, -9, -2, -11, -10, 12, 12, 16, -10, -15, 6, 4, -13, -12, 7, 0, -1, -1, 11, 6, 1, 11, -23, 2, -23, -17, 20, -2, 29, 1, 0, 22, -11, -6, 10, -1, 11, 15, 2, 17, 0, 13, -12, -12, 0, -4, 7, -14, -6, -23, 10, -13, 5, 21, 6, -2, -4, 2, -4, -1, -7, -17, 9, 22, 19, -5, -1, 2, 10, 5, -11, 17, -21, -6, -1, 5, 4, -15, -15, -17, 3, -1, 8, 5, -8, 12, 11, 6, 10, -1, -3, -21, 1, -6, -21, -7, 8, -12, -5, -19, 11, 16, 6, -7, -2, -23, -5, 0, -16, 13, 16, 12, 22, 2, 11, 4, 14, 3, -30, -3, -16, 1, -10, -12, 27, 0, -3, -23, 0, 9, 1, -4, -5, 8, 5, 31, 12, -8, 2, -17, -5, 9, -14, -8, -10, 12, -3, -9, 16, -4, -2, -8, 2, -12, -3, -8, -13, 6, 11, -5, 0, 8, 0, 22, 4, 11, -8, 6, -14, 5, 9, 6, 15, 2, -5, -2, 2, 9, -8, -6, 1, -1, -9, 10, 0, 3, 6, -14, -2, -6, 5, -2, 8, 8, 1, 4, 7, 15, 3, 5, -6, 1, 15, 15, -9, 9, 22, -2, -7, 13, 12, 22, 2, -6, -8, 8, 1, 9, 8, 7, 14, 8, -9, 8, 1, 8, -16, -9, -4),
    (-14, -5, 1, -19, -11, 32, -2, 1, -27, -12, -23, 0, -21, 6, 13, 1, -3, 11, -4, 11, 9, -24, -10, -6, -1, 0, -4, 15, -14, -9, -9, 2, 6, -20, 30, 6, 7, 7, -2, -9, -4, -15, 0, 5, 27, 3, -8, 13, 12, 11, -23, 11, -11, 18, 8, 1, -9, 5, -11, 0, -8, 13, 16, 2, 16, 13, 0, 7, 8, -28, 22, 9, 6, -12, -17, 12, -17, -11, 3, -7, 4, -19, -11, -1, 21, 12, -13, 7, -7, -20, -9, -4, 23, -9, -11, 12, -3, -7, -11, 6, -4, 4, 0, 2, 9, 3, -8, -17, -3, 17, 8, -6, 3, 8, -17, 13, 3, -18, 13, -9, -7, 12, -11, 9, -13, -19, 3, -8, 1, 3, 9, -6, 18, 5, -28, 12, 0, 0, -3, 0, 2, -10, -12, 16, 10, -8, -15, -20, 7, -16, 12, 4, 17, 4, -24, -22, 6, 28, 10, -14, -10, -3, -13, 8, -12, -16, 3, -5, 12, -8, -13, 10, -13, -2, -11, -11, 6, -8, 4, -8, 15, -4, -9, 0, -6, 0, -7, -13, 16, -9, -9, -5, -28, -10, -15, -7, -3, -3, -8, -7, 4, 4, -8, 6, -9, -10, 14, 5, 5, 3, 0, 4, -8, -8, 3, 11, 5, -33, -6, -4, -5, -14, -3, 8, -3, 1, 15, 9, 7, 12, -3, -6, -6, 9, -1, 15, -2, 11, -16, 13, -12, -8, -30, -10, -2, 5, -1, 11, 1, 7, -5, 1, -11, 11, 13, -4, 5, 0, -16, 13, 5, -6, 11, 9, -16, 8, -10, 10, -2, -16, -6, 0, 6, -7, -9, -3, 5, 14, 2, -2, 6, 0, -12, 11, 10, 0, -28, 5, 2, -18, -10, 6, -21, 16, 17, 23, -11, -6, -19, -9, 3, -1, 1, 3, -1, 10, -30, -2, 3, -15, 9, -4, -26, 12, 2, 18, 3, -21, 11, -16, 8, 1, 19, -7, 11, 14, -11, 2, 1, 16, -12, -12, 19, -3, -1, 3, 7, -23, -9, 4, 7, 2, -3, -3, -1, -11, -15, -24, 4, -1, 12, 10, -10, 8, -16, 13, -10, -3, -4, -18, -18, -1, 10, 11, 10, -19, -12, -15, 12, -1, 11, 10, 13, 13, -16, -3, -12, 17, -14, -18, 6, -6, 4, -3, 2, -20, -5, 2, 5, -18, 7, -6, -8, 5, -18, 1, 2, 12, -2, 14, 10, 9, -3, 17, -4, -10, 8, -9, -1, -14, -2, 2, -5, -12, 2, 3, -4, 3, 33, 2, 3, 21, -3, -6, -5, 7, -2, 10, 3, -11, -18, 14, -7, -9, -7, 10, -3, -3, 7, 11, -11, 11, -8, -12, -13, 13, -2, 7, -8, 1, -14, 9, -3, -6, -10, -7, -15, 10, -6, 21, -5, -14, 2, -9, 3, 6, 15, 7, -2, 11, -1, -10, 6, -2, 1, -2, 14, 1, -16, 4, 1, -4, -3, -6, -14, -1, 5, 7, -8, 8, -7, 1, -5, 5, 11, 3, -10, -2, -3, 6, 6, -7, 3, -6, -6, 9, -1, 19, -4, -21, -4, -5, -1, -5, 15, -8, 5, 17, 7, 2, 9, 6, 10, 5, 7, 0, -1, 9, 3, 0, -12, 11, 3, -5, 13, 4, -9, 0, -2, -10, 3, 2, -7, 11, -9, 6, -9, 5, -3, -14, 1, -11, -11, -8, 0, 12, -11, -19, -11, -5, 0, -12, 8, -6, 15, 6, -5, -6, 4, 1, -6, -7, 18, -16, 1, 9, -19, -23, 5, 9, 4, 13, -3, -3, -7, 19, -9, 0, -7, 23, -6, 11, -5, 6, 10, 12, 6, 4, 0, -4, 2, -3, 6, -1, -13, -10, -11, -2, 6, -16, 23, 19, 10, 5, 4, 12, -10, 3, 5, -6, 4, -14, -12, -6, -2, -7, 1, 6, -3, 5, 4, 10, -15, -5, -6, -5, 2, 18, 0, 2, -2, 11, 1, 19, 9, -8, 0, 13, 0, 13, -2, -4, -12, -8, -18, 10, 23, -19, 12, 5, 8, 16, 8, 2, 6, 1, 10, -5, 17, -19, -6, -7, -2, 3, 0, 8, -13, 7, 1, 0, -14, 3, -6, -2, -1, 11, 13, -3, 9, 2, 1, 12, 14, -6, -5, 8, -10, -10, -4, 12, -16, -13, -4, 2, 17, -17, -5, -2, -13, 9, 16, -5, 4, -2, -1, 16, 13, -11, 0, -5, 9, -4, -10, 21, -14, 0, 11, 8, -16, -8, -3, 6, 8, 1, 5, -1, -11, 2, -9, 6, 3, 2, -2, -3, -3, 3, -7, 1, -12, -9, -16, 5, 6, -24, -14, -25, 3, 13, 3, -4, 9, -1, -9, 5, -6, 8, -7, 14, -2),
    (-14, 5, -14, 2, -10, -14, 11, -13, -29, 10, -9, 20, 11, 12, 6, -6, -5, 20, 9, 13, 14, -20, 8, 4, -3, -7, 0, 8, -4, 8, 8, -21, -9, -2, -13, 9, -8, -4, -6, 14, -1, 8, 3, -12, 13, 2, -9, -3, -7, 25, 0, 4, -8, -9, 5, 14, 0, 7, -2, -8, 4, -21, -23, -28, -18, 5, 18, 1, 24, -15, -27, 2, 19, -4, -14, -4, -3, -14, -2, -7, 1, 10, -14, 1, -32, -6, 5, 14, 0, 39, 5, 2, -2, -7, -7, -4, -16, 25, 3, 11, -5, -2, 3, 10, 21, 8, -2, -3, -5, -26, -19, -16, 11, 7, 0, -2, 17, -36, -22, 13, 10, 5, -18, -18, 10, -19, -5, -24, -3, 8, -5, -2, -9, -3, 18, -1, 3, 26, 2, -7, 2, 12, -4, 9, -24, 21, 20, 9, -16, -5, -11, 15, 20, 8, 17, 12, 7, -24, -5, -4, 2, 11, 10, -27, 12, -14, -2, 7, 10, 6, -32, -15, -10, -12, -14, -20, -20, -1, -5, -2, 7, 9, 20, 7, -3, -2, 11, -7, 8, 4, 0, 18, -42, 10, 8, -5, -9, -35, 16, -9, -22, 7, -12, 16, 18, -6, -1, 7, -17, -1, -2, 16, 18, -18, 2, 15, 8, -16, 1, -9, -11, 11, -10, -6, -3, 1, -44, 1, -12, -14, -6, 24, -11, 6, 1, -2, -14, 9, -8, 3, -27, 10, 18, -11, -22, -29, 1, 0, -4, 25, -13, 9, 4, 5, -6, 1, 0, 16, 17, 15, 17, -31, -36, 6, 15, -23, -8, -4, -14, -25, -1, 5, -2, -6, -13, -3, -10, -5, 1, 26, -10, 10, 9, -21, 6, 22, 2, 1, -14, 19, 7, 5, -29, -20, 2, 23, 9, 17, -12, -3, -1, -3, -3, -5, 0, 19, 16, 5, 4, -6, -19, 18, 7, 2, -23, -9, 3, 3, 1, -1, -20, -3, 6, 2, 7, -3, -6, 15, 13, -2, -1, 3, 0, 3, -3, -8, -29, 22, 7, 12, -25, -9, -1, 19, 0, 23, 11, -5, -6, 1, -16, 17, 1, 17, 4, 8, -8, -18, -10, 8, 1, 10, -24, -7, 2, -1, -1, 9, -26, -11, 7, 15, -3, 3, -1, 3, 0, -1, 0, 0, 3, -2, 3, -6, -30, 12, 6, -21, -7, -67, 5, -9, -1, 2, -17, -8, -1, -4, -7, 11, 10, 15, -6, -6, 10, -40, -20, 12, 3, 1, -14, 0, -7, -17, 13, 10, 13, -11, -46, -2, 9, -12, -8, 7, -10, 22, 15, 3, -6, 28, 10, -10, -7, 14, 2, -9, -17, -42, 10, 11, -3, 16, -33, 2, -3, 7, -20, 0, 13, 8, -2, 6, 6, -36, -29, 18, 16, -29, -17, 11, -1, -5, 13, 2, -5, -1, -10, -3, 0, -14, -18, 23, -16, -7, 21, -14, 4, -2, 7, -9, 8, 7, 9, -2, -20, -23, 6, 8, -6, 8, -7, -10, 18, -6, -2, 1, 21, 7, 17, 5, -4, 10, -26, 11, 18, -9, -19, -7, 1, 14, 13, -4, -16, 5, -3, 5, 0, -23, -1, 8, -11, 11, 8, -25, -2, -5, 2, 13, -9, -2, -1, 27, -22, -10, 5, 15, -2, 13, -9, 5, 10, -9, 13, 10, -1, 14, 10, 1, -2, 5, -12, 0, 11, 7, -18, -7, 1, -4, 8, -5, -8, -6, -2, 7, 7, -9, 10, 15, 7, 4, 7, 11, -4, -14, -19, -10, -9, -2, -4, -21, 4, -1, 1, 4, 10, 4, -16, 6, 8, -15, -7, 3, 9, 16, -15, -18, 4, -19, 5, 10, 12, -12, -23, -12, 2, -8, 11, -5, -9, 1, -38, -22, 11, 7, -17, 0, 10, -1, -3, 2, -16, -10, -1, -3, -8, 14, 9, -29, 1, 4, 6, 13, 7, 5, -10, -4, 10, -8, -20, 7, 10, 10, -25, 2, -10, -28, -8, -5, 6, -37, -8, -26, -1, 3, 17, 8, -9, 8, -43, -4, -8, -13, -33, 2, 0, 12, -6, -4, 18, -10, 4, -3, -12, 13, 9, -5, -10, 1, 7, 2, -11, 8, -19, -6, 18, -4, -9, 5, 22, 5, -5, -3, -7, -16, -9, -14, -7, -5, -22, -15, -9, -11, 4, -9, -12, -3, -23, 5, 1, -2, -19, -9, -2, -1, 9, -13, 17, -2, -7, 4, -9, 8, 9, -12, 6, -7, -5, -22, -5, -6, 11, 6, 9, -17, 16, -16, 16, -6, 4, 19, -11, 2, -11, 5, 10, 6, 4, 0, 6, -4, -7, 2, -17, -9, -6, 10, 1, -7, -21, 6, -8, 11, 18, -4, 7, -11, -22, 0, 2),
    (12, -6, -1, -5, -19, -12, 3, -6, 1, -1, 25, 4, 22, 14, 8, -2, -2, 5, -31, -8, 16, -3, -10, 3, -10, 6, 13, -6, 19, -13, 6, 7, 7, 14, 0, 3, -31, 0, 8, -7, 8, 1, 0, 9, -18, -4, 5, -8, 3, -11, -9, 15, -50, -2, -3, 15, 10, 12, 13, 1, 21, -3, 9, 11, -5, -2, -30, 3, 11, 12, -17, 18, -12, 5, 13, 15, 5, 1, -7, 10, 8, 12, 9, 1, -9, 9, -13, -52, -4, -14, -2, -4, -16, 1, -16, 0, 6, -20, -8, 16, -7, 15, -10, 16, -8, 18, 18, 23, 5, 3, 11, 18, -27, -9, -34, 5, -5, 14, -1, 0, -7, -10, 10, 4, 2, 8, 2, -22, 0, 15, -11, -2, -3, 13, -6, -67, 5, -13, -7, 4, -4, 12, -32, 1, 5, -3, -4, 24, -12, 27, -13, -23, -9, -7, 12, 22, 13, -31, 0, -8, -34, -8, -27, -14, 22, 7, -3, -20, -21, 7, 3, 2, -3, -9, 3, 1, -1, 13, -1, -11, -12, 5, 17, -30, 18, 26, -15, 10, 1, -9, -23, 6, 4, -16, 9, 8, -10, -33, -10, -5, 12, -15, -4, 4, 5, 9, -10, 14, -3, 8, -25, -1, 1, 7, -2, 7, 5, -3, -3, -1, 3, 7, 1, 1, -14, 17, -7, 11, -12, -8, 4, -28, 10, 11, -7, 7, 20, -6, -4, 4, 16, -14, 4, 19, -25, 4, -13, 10, 0, -14, 11, 2, 18, 15, 3, 8, 4, -4, -2, -8, 8, 5, -9, -10, 0, -10, -2, -2, -3, -28, 10, 3, -15, 7, -4, 2, 5, 10, 0, -51, -11, -12, 7, 6, 20, 0, -9, -4, 6, -13, 0, 13, -24, -5, -8, -11, -4, -17, 20, 14, 3, 3, 11, 21, 14, -13, -1, -12, 7, 3, -8, -9, -12, -7, -13, -7, -6, -21, -6, 23, -15, 4, 3, 15, -4, 5, -7, -47, -10, -18, 10, 9, 19, 3, -31, -13, 12, -10, 8, 21, -17, -4, -20, 2, 4, -12, 14, 24, 5, 2, 7, 0, 18, 5, -24, 6, -4, -6, -8, -5, -18, -12, -27, -23, -7, -18, -6, 27, -13, 11, -3, -1, 9, -14, -29, -18, -7, 15, 1, 12, 12, -9, -21, -9, -4, -16, -10, 6, -7, -8, 8, 9, -6, -11, 1, -10, 5, 3, -7, -8, 6, -8, -4, -12, -4, -9, 1, -3, 0, -4, -7, 24, -8, -10, 4, 10, -3, -2, 4, -4, 1, 17, 6, -24, 2, 2, -9, 22, 14, -4, -26, 11, 12, -19, -9, 18, -17, -3, 1, 3, -17, -31, -7, 9, 8, -4, 11, -6, -2, -2, 2, 2, 4, -8, -4, -1, 6, 1, -2, -7, -3, -10, -8, 12, -10, -5, 3, 1, 7, 19, -11, -28, -13, -10, -1, 1, 22, 5, -19, 9, 12, -8, -4, 11, -35, -8, 7, -4, -1, -23, 11, 3, 10, 2, 16, 9, -2, -11, -14, 10, 7, 2, -5, -10, -10, 7, -6, -25, -10, -17, -15, -5, 0, -6, -12, 11, -2, -7, 2, -27, -21, -11, 3, 11, 19, 14, -9, 0, 13, -12, -17, -3, -10, -16, -5, 15, 4, -28, 7, -13, -9, 14, 13, 2, -2, 2, -6, 6, 6, -3, 2, 12, -12, 3, -8, -6, -1, -9, -16, 12, -6, 8, -13, 8, -9, -12, -5, -18, -26, 0, -1, 21, 7, 8, -5, 0, -18, -4, -3, 14, -11, -9, 5, 14, -17, -12, 2, 7, 10, 6, -3, 7, -12, 5, 13, -24, 14, -7, -4, 3, 3, -23, -3, 5, 6, -2, 6, -2, 6, -17, 2, 17, -4, 8, 15, 12, 8, 5, 3, 5, 5, -12, -10, 14, -2, -8, 9, 14, -17, -5, -2, -6, -12, -23, -2, 8, 8, 6, 9, 1, -11, -1, -5, 3, 7, 5, -10, -2, 3, -17, 11, -7, 8, -6, -4, -1, 1, -17, 16, 0, 13, 7, 3, -9, -10, 7, -5, 1, 22, 0, -19, 5, 4, 2, -4, -3, -10, 10, 0, -6, -17, -9, -3, -2, 5, 19, 17, 4, -2, 8, -8, -1, 10, 0, 7, -6, -7, -5, 9, 8, -2, -18, -11, -1, -1, -7, 7, 14, -6, 4, 3, -6, -5, -2, 11, -6, 18, -15, 8, 2, -2, 0, 0, 5, -16, 4, 12, 11, -7, -6, 0, -8, 4, 7, 6, 1, -8, -15, -6, 8, 8, -7, 5, -1, -7, 11, -10, 7, -5, -8, -16, 10, -10, -15, -5, 3, 3, 2, -5, -6, -23, -2, 6, 4, 4, -8, -1, -12, 0),
    (-6, 17, 0, -14, 4, -25, -10, 22, 34, -13, 9, -9, 15, 13, -14, 20, -7, -1, -26, 34, -28, -15, 19, 4, -2, 21, 6, -5, 2, -4, 4, -6, 9, -2, 5, -16, -18, -31, 0, -17, -1, 18, 9, 0, 4, -10, 25, -27, 0, 3, -3, -23, -9, -36, 1, 25, 28, -2, 11, 6, 4, -14, -10, -2, -16, 4, -18, 10, 3, -20, -18, -7, -7, -5, -7, -12, 14, -11, -16, -17, 0, -8, -11, 9, -12, -9, 3, -25, -3, 13, 15, -8, -2, -11, 25, -2, -4, -19, 0, -21, -4, -13, -8, 10, 10, 4, 2, 18, -12, -30, -9, -17, -4, -16, -13, -5, 9, 0, -22, -14, -13, -8, -9, -8, 7, -37, -8, -16, -5, -5, -35, 1, -15, 7, 10, -31, -5, -3, 19, 15, -2, -2, 11, -16, -10, -35, 2, -6, 4, -4, -10, 16, 3, 0, -1, 10, 4, -21, -23, -20, -19, -26, -8, 6, 18, 8, -10, -17, -5, -15, -10, -13, -17, -14, -19, -5, -15, -7, -2, 6, -18, -5, 0, -32, -10, 5, 24, -3, -10, -8, -10, -13, 10, 0, -2, 0, -10, -10, -1, 8, 14, 22, 16, -2, -5, 13, 2, -2, -13, 3, -24, 20, -6, 15, -4, -3, -5, -21, 3, -18, 8, -5, 19, -19, 24, 10, 6, -1, -6, -16, -10, 9, 13, 11, 10, -9, -25, -13, 11, -5, 13, -19, 10, 10, -16, -32, 3, 15, 19, 19, 11, 4, -3, 5, 3, 1, -24, -9, -15, 3, -13, 6, -2, -2, -3, -22, 0, -18, 15, -16, 10, -5, -4, 19, -7, -2, -27, -12, -32, -8, 7, 8, 14, -1, -17, -5, -4, -7, 9, -17, 1, -1, -5, -2, -16, 16, 6, 5, 7, -16, -15, -12, 10, -14, 17, -14, -17, 6, 3, 0, -17, -16, -9, -12, -6, -17, 13, -30, -2, 2, -8, 12, -11, 12, -5, -14, -41, -5, 20, -1, 14, 3, -6, 12, -7, 4, 12, -10, -11, 1, -8, -15, -1, -2, -3, 14, 5, 2, -1, 3, 19, -2, 3, -37, -7, -5, 14, -10, -4, -18, 10, -12, -6, -25, 5, -20, 9, -11, -9, 17, -22, 17, -5, -20, -39, -27, 22, 8, 15, -3, -2, -10, 1, -10, 9, 9, -3, 12, -5, -16, 8, -1, 10, 20, 12, -5, 5, 7, 2, -14, -14, -6, -10, 19, -1, 10, -3, 2, 10, -7, -8, -17, 3, 1, 12, -8, -12, 12, -5, 0, -17, 3, -19, -4, 23, 8, 4, -12, -11, -11, -3, 5, 19, -8, -4, 12, -25, -23, -9, 10, 17, 21, 1, 6, -21, -3, 4, -4, -1, -11, -12, -4, -9, -7, 8, -9, 7, -14, 1, -19, 4, -17, 3, 9, 0, 20, 15, 12, -10, -17, -26, 5, 17, -5, -2, -20, -29, -17, -18, 11, 14, -1, 3, 1, -16, -17, -11, 16, 10, 17, 3, -19, -15, 10, -1, -9, 3, -6, -8, 8, 3, 7, -14, -23, 12, -10, -14, 0, 0, -24, 9, -3, -1, 1, -8, -3, -12, -15, -28, 4, 12, 7, 5, -8, -15, -2, -11, -9, 8, 27, -9, -1, -9, 2, 3, 8, -11, 20, 5, 2, -8, 1, 7, -19, -7, -8, -14, -4, 14, -7, 7, -8, 3, -18, 5, 4, 13, -10, -2, 7, -19, 7, -7, 3, -16, -19, -12, 1, 20, -1, 1, 2, -6, -20, -11, -5, 21, 6, -5, 10, -3, 2, -11, -14, -3, -3, 18, -2, -9, 12, -2, -21, 1, 11, -12, -4, 6, 1, -1, -7, 7, -5, 2, -16, -3, -8, 6, -1, -3, 1, -8, 7, -5, -10, -16, -15, 20, 3, 3, -10, -13, -3, -2, -1, 10, 6, -3, 10, -1, -16, 1, -15, 10, 18, 14, -11, -28, 13, -7, -23, -10, -3, 4, -4, 6, -6, 7, 8, -4, -3, 6, -8, -4, -8, 18, -17, -10, 12, -16, -5, -13, -5, -30, -15, 4, -5, -2, -19, -8, -8, -18, 9, 10, 11, 10, -10, 4, -27, -18, -10, -17, 16, 8, 3, -12, 8, 5, -12, 8, -5, -6, -1, -6, -8, 10, 1, -14, -3, -5, 0, -1, 1, 17, -8, 6, -9, -17, -3, -22, -8, -2, -1, 10, 5, 7, -14, -12, 2, -24, 1, 15, 17, 3, -32, -6, -25, -17, -8, -25, 5, 8, -11, 3, 7, -6, -8, -13, -13, -11, 5, -9, 3, -8, -3, 12, -2, -27, 4, -7, 3, 10, 6, -10, 7, -19, 6, -15, -3, -19, -8, 11, 4, 14, -4, -8, -11, -21, 0, -11),
    (6, -1, 2, 11, -1, 9, 2, -19, -34, -5, 0, 12, -13, 5, -8, -4, -16, 4, 1, -2, 19, 13, 12, 1, -23, -2, 16, 5, -10, 11, -11, -8, -16, 5, -7, -1, 7, -6, -18, 9, -12, -20, 11, 3, 8, 1, -11, -8, -5, -13, 22, 13, 16, 3, -6, -27, -14, 9, -20, 10, 6, 13, -2, -6, -26, 4, 9, 1, 26, 10, 17, 7, -35, -1, 2, -1, -6, 19, 9, 20, 17, 1, 17, -13, -21, 4, -6, 6, -1, -4, -6, 27, 9, -12, -6, -8, -15, 10, 3, 8, 16, 12, 3, 3, -26, 11, -21, -33, 8, 7, 5, 11, -4, -9, 3, -6, -3, 4, 13, 9, -19, -9, 5, -2, 11, 17, 2, 47, 9, -11, 1, 2, -4, -6, -8, 10, 13, -11, -28, 7, 8, 1, 13, -4, -20, 9, -6, 7, -3, 0, -2, -10, 2, 21, -20, -13, 11, 17, -3, -1, 4, -13, 1, -20, -9, -5, 5, 4, -9, -4, 2, 0, 7, -6, 19, 4, 12, -11, 6, 2, 1, 0, -22, 9, 10, -15, -6, -15, -3, 0, 7, -12, 27, -11, -12, -14, 4, -3, -3, -9, -7, -9, -30, -18, 16, -11, 14, 3, 18, -7, 4, 5, 4, -12, -9, 6, -24, 15, 15, 9, -1, 20, 1, 6, -7, -22, -11, -7, 26, 4, -20, 4, -20, -1, 4, 0, -4, -19, 26, -28, 2, 12, -12, -27, 22, 10, -4, -3, -17, 16, 0, -1, 17, 10, 2, -7, 27, -7, 13, -15, 2, -25, -10, 9, -33, -2, 18, -2, -26, 11, 5, 19, 10, -31, -13, -5, 9, 13, -1, 5, -11, -16, 1, -17, -6, -28, 37, -17, -6, -3, -7, -19, 10, 6, -19, -14, -3, 27, -5, -15, 12, 8, 3, -1, 32, 10, 10, -17, 0, -33, 2, 9, -17, -4, 6, -19, -8, 5, 11, 17, 6, -28, 5, -15, 13, -3, 15, 6, -14, -6, 2, -15, -12, -34, 10, 4, -7, -6, -6, -28, -2, -3, -2, -8, -8, 3, 4, -16, 12, 11, -8, 4, 23, 16, 6, -7, -21, -4, 10, 10, -20, 3, 0, -17, -12, 6, 2, 1, 10, -28, -9, -17, 12, 5, 8, 26, -37, -16, 13, -4, -4, 14, 14, 3, 21, -8, 0, -22, 2, 0, -31, -18, 6, -26, -22, -8, 0, -1, -18, 10, 9, -12, 5, 2, -5, -5, 10, 18, -24, 9, 10, -19, 4, 9, 6, -3, 8, -31, -3, 0, 20, -11, -16, 13, -38, -6, 9, -15, -4, 5, 22, -44, -7, 16, -12, -22, 22, -4, -37, -17, 1, -8, 3, 8, 22, -11, -23, -1, 4, -11, 19, -6, 0, -32, 1, 25, -27, -5, -3, -11, -28, 7, 24, 4, 16, -31, -15, -16, 15, -7, -2, -14, -7, -21, 22, -11, 8, -8, 23, -22, -3, 6, 6, -12, 29, -6, -29, 7, -1, -8, 7, 7, 22, -19, -16, -16, 19, -9, 13, -22, 0, -4, 1, 31, -9, -9, -9, -7, -23, 10, 13, -13, 13, -28, 1, -20, 17, 3, 19, -4, -10, -23, -1, -12, -12, -15, 21, -12, -3, -15, 13, -23, 3, 7, -8, -9, 11, -7, 4, 11, 19, -14, -16, -6, 21, 15, 10, -9, -1, 3, 10, 19, -17, -7, 16, -16, -36, 17, -19, -13, 9, -27, 9, -7, -1, -6, 12, 18, -12, -19, 2, -20, -6, 4, 0, -19, -2, -25, -2, -18, 1, 11, -1, 3, 21, 3, -32, -2, 9, -41, -19, 12, -2, -50, 13, 13, -20, -7, -9, 14, -1, 3, -19, 6, -12, 4, -1, -24, -6, -5, 21, -49, 13, -15, -8, 13, -14, -23, -1, 1, -6, 8, -1, -15, -22, -12, 6, -46, -14, 8, -6, 11, 11, -11, -16, 1, 16, -33, -24, 17, -6, -35, 15, -5, -20, -5, -13, 10, -4, 6, -8, 3, -31, 15, -12, -21, 4, 10, 13, -30, 18, 3, 12, 2, -17, -27, 4, 1, -11, -3, 15, -10, 2, -10, 5, -17, -13, 11, -24, -4, 17, -7, 18, 12, 13, -17, -34, 2, -12, -28, 9, -9, 13, 3, 11, 9, 13, 6, -7, -2, -17, -17, -4, -18, 7, 20, -13, -22, 12, 9, 13, 9, 9, -8, 0, -5, -13, -5, 2, -7, 6, -5, -1, 6, 2, 17, -4, 12, 14, -12, 0, 1, 11, -13, -31, 18, 1, -4, 13, -5, 17, 3, 10, -10, -2, -1, 2, -14, -4, 2, -7, -24, 11, 9, -4, 0, 10, 0, 6, -1, -7, -10, -5, -7, -3, 21, 17, 12, 4),
    (-17, -5, 5, -3, 13, -5, 11, -11, -19, 1, -19, 2, -17, 2, -8, -20, 7, 15, 13, -8, -9, 6, -4, -12, 3, -19, 13, -5, 13, 0, 4, 1, -7, -7, -10, 11, -7, -4, 17, -15, 12, 8, 6, -13, 5, 11, -15, 9, 17, 0, -10, -2, 5, -14, 20, -7, -18, 2, -12, 3, -19, -4, -7, 6, 5, -1, -2, -9, 8, 5, -7, -7, 30, 1, 20, -11, -1, -20, 4, 2, 3, -9, -16, -1, 19, 0, 7, -11, 4, 20, 4, -19, 12, 18, -8, 8, 9, 12, 7, -8, 21, -14, 17, -12, -20, -12, 4, -6, -14, 10, 4, -11, 6, -4, -13, 7, 17, 1, 1, -16, 9, 19, 9, -16, 3, -9, -2, -2, -1, -7, 2, -8, 1, 1, -6, 6, -5, 23, 8, -9, 4, 9, -11, 24, 19, 6, -1, 2, -1, -8, 12, -4, -6, -11, -12, 0, 1, 0, 6, -3, 3, -4, 2, 6, 12, 9, 0, 7, 5, 11, 12, -13, 16, 9, 9, 9, 12, -19, -11, -11, 3, -4, -4, 1, -5, -3, 8, -3, 12, 1, -9, 20, 15, 12, 7, 4, 0, 8, 5, -14, -17, -33, 13, 5, -32, 2, 6, -24, 2, 16, 7, -12, 0, 6, -6, 10, 8, 6, 15, -9, 8, 16, 5, -3, -28, -21, -8, -13, 5, -2, 11, -41, 9, 16, -17, 8, 11, 1, 9, 3, 16, 7, -13, 9, -1, 1, 16, -20, -11, -10, 3, -1, -25, -9, -3, -9, 1, -10, -16, 6, -13, -1, 3, 0, 18, 35, 17, 1, -2, -14, -3, -12, -2, -23, -10, -18, 11, 4, 12, -12, 4, 8, -5, 5, 0, 0, 0, 8, 8, 4, 2, 1, 36, 0, 6, -15, -11, -8, -11, 11, -1, 8, -10, -17, -5, -8, -12, -5, 11, 6, -5, -2, 10, 20, 18, 8, -5, -4, -14, -24, 9, -4, -5, -6, -2, 6, -4, -15, 1, 1, 6, -11, -3, -8, -5, 12, 13, 12, 0, -4, 14, -4, 16, -12, -8, 6, -17, -2, 5, -7, 2, -19, 2, -10, -10, 4, -5, 4, -9, -8, 16, 16, 11, 15, 4, -7, 13, -8, 0, -9, 3, 1, 9, -3, -1, -16, -5, 18, 11, -10, -5, -14, 12, 6, 1, 20, 3, 2, -2, 18, 13, 8, 4, -14, 7, -2, -8, -9, 11, -23, -8, -2, 2, -12, -10, 21, -8, -3, 7, 11, 9, -1, 1, 3, -12, 5, -18, -20, -23, -23, -12, -23, 12, -29, -5, 11, -23, 15, -1, 12, 12, 8, 20, 7, -5, 13, -14, -8, 13, -21, -13, -11, 7, 10, -9, -1, 14, -16, -9, -9, 20, 4, -2, -4, 1, -12, 12, 22, 19, 7, 17, -28, -24, -2, -7, -32, -4, -9, -6, -21, 0, -40, -16, 2, -9, 16, -12, 11, -7, 15, 16, -10, -11, 2, 27, -18, 5, -29, 5, -4, -9, 8, -3, 4, 8, 7, -4, -20, 5, 8, 4, 8, -12, -12, 7, 25, 10, 11, 8, -27, -18, -22, 0, -9, -4, -1, 2, -14, -5, -35, -9, 7, 0, 17, 9, 10, 4, 15, 14, -11, -6, -11, 7, -12, 7, -9, 7, 4, -2, 5, -9, 4, 10, -1, -1, 7, -2, 11, -10, 5, -11, -7, 7, 14, 4, 19, 3, -6, 2, 2, 5, -20, -4, -5, -10, -14, 9, -7, -5, 0, -14, -4, -1, -13, 14, 7, 16, 30, 3, 6, -11, -5, 4, -1, -13, -12, 12, -5, -2, -5, 15, -18, -5, -12, -24, -18, 0, 20, -9, -13, -3, -4, 9, 15, 7, -5, 7, -12, -16, -1, -26, 3, -5, -19, 18, -14, -20, 15, 7, 9, -4, 5, 7, 19, 14, -1, 1, 12, -21, -18, 8, -7, -11, 7, 1, -14, -19, 2, 12, -13, -1, -22, -17, -15, 10, 5, -13, -27, 8, 17, 10, 26, 14, -17, -4, -11, -20, -13, 9, 10, -6, -12, 9, -10, -31, 20, -8, 8, 0, 9, -6, 11, 21, -6, -15, 2, -12, -11, 7, -7, -10, -3, -6, 2, -8, -8, 25, 8, -17, -27, 2, 2, -7, 3, -17, -8, 9, 13, 1, 8, 23, 11, -4, -19, 2, -8, 9, 5, -16, 1, -10, -18, -17, 8, 6, 24, 4, -4, -11, 4, 21, -3, -12, -17, 4, -15, 2, -8, -18, -8, 4, -4, -9, 1, 11, 9, -16, -7, -6, 12, -3, -10, 5, 0, -9, -1, 2, 10, 11, -9, -33, -26, -1, -33, 20, 4, -18, -4, -6, -16, -21, 2, -7, 6, -6, -2, 14, -5, -3),
    (1, -6, -7, 7, 0, 6, 13, 1, -15, 2, 3, 13, -25, 12, -7, 1, 7, -12, -3, -18, 9, 15, 2, -25, 4, -36, 17, -4, 20, 0, 8, 4, 22, -7, 2, 2, -14, 3, 13, 1, 13, -2, 12, -9, -31, 11, -20, -2, -13, -19, 18, 3, 9, 2, -7, -6, -16, 11, 0, 3, -30, -6, 13, 27, -35, -8, -8, -1, -12, 1, -13, -25, 20, -25, 16, -32, 8, 3, 3, 17, -1, -8, 16, -3, -13, -12, 5, -13, 2, -1, 12, -25, -4, 3, -6, -2, -8, -12, 14, -6, -26, -18, 2, -31, -39, -10, 5, 2, 2, -4, -3, 12, -24, -8, -12, 4, -7, 16, 9, -13, 11, -20, 18, -16, 12, 23, 3, 2, -1, -6, 10, 15, -1, -8, -3, 0, -1, -4, -3, -20, 12, 6, 15, 2, 5, -23, -1, 0, -6, -11, 5, -21, -31, -13, -7, -17, 1, -4, 9, 25, 11, -9, 4, 3, -7, 6, -2, 1, -4, -10, 15, -17, 22, 9, 18, -2, 3, -6, 16, 13, 4, -11, -21, 4, -2, -8, -15, -10, 10, -15, 0, -3, -10, 9, 18, -10, 12, -16, -4, 4, -8, -5, -16, -3, 1, 1, -2, 15, -3, -8, -14, -7, 4, -8, 31, -31, 6, 0, -9, -1, -2, -16, 20, 2, 25, -32, -27, 2, 8, -11, -4, 1, -13, -3, 7, 5, 5, -4, -19, 4, -9, 9, 27, -14, 11, -22, -10, 3, 10, -4, -10, -2, -29, -7, -12, 13, -6, -13, -11, -7, 24, -4, 6, -39, 19, -24, -14, -11, -1, 3, 16, 14, 7, -25, -32, 11, 8, -1, 3, 5, -17, -7, 24, -5, -3, -19, -12, 4, 6, 7, 7, -20, -24, -20, 5, -29, -2, -5, 1, 7, 1, 6, -13, 2, -9, -16, -12, -5, 27, 30, 12, -17, 24, -27, 1, -14, 11, 13, 13, 4, 3, -3, -9, 9, 12, -7, -8, 2, -12, -6, 16, -6, -16, -20, 7, 14, 11, 12, -5, -35, -17, 0, -8, -24, 3, -20, 10, 10, 1, 8, 6, 8, -10, -6, -16, -6, 23, 13, 16, -8, 26, -15, -3, -12, 11, 13, 11, -2, 6, 7, -21, -2, -1, -10, 3, 9, -20, -9, 5, -7, -5, 2, 6, 20, -29, 13, 22, -24, 6, -47, 15, 13, 28, 1, -14, -9, -2, 6, -4, 19, 10, 14, -11, -10, 4, -37, 25, 8, 11, -4, -12, -11, 9, -6, 33, 7, 12, -25, -57, 9, -11, -10, -3, -1, -13, 0, -8, 8, -2, 7, 0, -7, -6, 5, 14, -15, -9, -18, 3, 23, 18, 14, -20, 12, -10, -17, -12, 14, 11, -3, -34, 2, -1, -13, 19, 0, 14, -31, -17, -8, 12, 11, 19, 5, 12, -19, -49, -19, 19, -14, -12, 27, -17, 3, 24, 3, 7, -13, -5, -1, -12, 14, -4, -25, -6, -25, -5, 12, 0, -15, -20, 6, 1, -5, 3, 14, 7, -16, -22, -5, 14, 26, 8, 1, 18, -42, -14, 0, 7, 13, 15, -2, 2, -14, -26, 2, 19, -21, -7, 25, -11, -7, 9, -14, 0, -11, -4, 9, 0, 14, -14, -36, 2, -2, 4, -5, 8, -6, 2, 10, -7, -4, -8, 15, 3, -10, -1, -3, 16, 12, 13, 9, 6, -3, -9, -1, 4, 2, 9, -10, -5, -3, -6, 15, 1, 1, 3, 10, -7, -10, 9, -18, -9, 6, -6, 20, -12, -11, 8, -20, -10, -28, -4, 9, 14, -4, -14, -15, 7, -3, 0, 7, 2, 16, 0, -4, 0, -13, 1, 15, 8, -17, -19, -21, -1, 3, -1, -7, 19, -6, -11, -26, 14, -11, 3, 7, 8, -15, -8, 14, -7, -4, 7, -12, -7, 9, 2, -34, -13, -21, -1, 11, 3, 0, -23, 3, -3, -17, -4, 28, 14, -5, 0, -3, -1, 7, 0, -8, 11, -3, -7, -26, -13, 19, -9, 6, 16, 8, -23, -1, 8, -22, 3, 2, -10, -2, 8, 8, 8, 5, 10, 3, -12, 21, 11, -30, -5, -7, -6, 14, 4, 2, -18, 15, 15, -17, -18, 22, 4, -1, -2, -3, -1, 13, 11, -6, 16, -17, -10, 0, 8, -9, -5, 4, 12, 7, -25, -7, 11, -4, -8, 4, 12, 8, -1, -11, -1, -6, -7, -2, -14, 15, 4, -22, 10, 3, -8, 17, -4, -12, -8, 3, 12, -12, -22, 15, 9, -1, -4, -13, -5, 6, 8, -3, 17, 8, -11, -9, -4, -4, 2, -2, 4, 6, -22, 13, 4, -1, -17, 15, -16, 0, -3, -2, 1, -9, -5, 11, -3),
    (6, -26, 5, 8, 12, 4, -16, 23, -20, 5, 0, 6, 2, 4, -5, 20, 11, -13, 17, -10, -7, 13, 11, -1, -14, 8, -9, -14, 12, 11, 18, -1, 2, 9, 19, 3, -13, -17, 8, 15, 8, 6, 8, -13, -1, -10, -3, -22, -8, -25, 1, -9, 5, 18, 0, 8, 7, -10, -5, 5, -7, 7, -18, -4, 20, -11, 10, -6, -40, 1, 12, -6, -19, 6, 4, -24, 13, 15, -1, 2, 1, 4, 15, 1, -23, -20, 23, 7, -4, 7, -6, 2, -5, -17, -15, 4, -4, -6, 5, -3, -40, -4, -9, -13, -9, 1, 7, -13, 9, 8, 1, 3, 25, 1, -5, -3, -31, 3, 9, -7, 2, 12, 17, -5, 16, 14, 12, 9, -11, 9, 8, 6, -27, -19, -3, 19, -2, -29, 0, 15, 10, -4, -3, -8, 7, -6, 3, -1, -17, -11, -18, -1, 13, -3, -7, -21, 7, 5, -1, 9, -8, -13, 11, -2, -33, 18, 4, -7, 10, 11, 3, 10, 6, 7, 14, 18, -4, 16, 10, -1, -6, 8, -15, 2, 7, -2, 4, 5, 10, 1, -4, -6, 7, -9, -15, 10, 12, 18, -15, 14, -8, -9, 14, 7, 5, 12, -4, -14, -7, -19, 7, 3, -9, 23, 0, -18, 7, -14, 9, -3, -10, -17, 15, -12, 4, -7, 26, -8, -17, -24, -8, 5, 10, -14, 1, -31, 5, -24, 10, -9, -17, -26, -10, -9, -4, 5, -1, 12, 5, 6, 4, 4, 15, 4, -3, -22, -7, -14, 5, -2, -10, 4, 13, -28, 2, 12, 8, -14, 10, 13, 4, -10, -2, 14, 22, 10, -23, -13, -13, 0, -3, -7, -8, -11, -4, -40, -26, -14, 8, -21, 1, -24, -3, 3, -10, 0, 1, -4, 28, -4, 1, 2, -13, -9, 1, -6, -24, -1, -11, -3, 0, -24, 5, 12, 0, -11, -2, 14, 0, 13, 2, -9, 5, -3, -26, -19, -3, 7, 0, -5, 1, -2, -21, -15, 5, -7, 0, -13, 15, -24, 7, 8, 1, 3, -8, -13, 7, -17, 9, 1, 2, -5, 7, -33, -5, -1, -22, -1, 15, -11, -5, 21, -15, -25, 11, 17, -6, -11, 9, 6, 18, 10, -13, 18, 4, -6, -7, -13, 13, -8, 2, -5, 2, -22, -5, -11, 6, 13, 4, 22, 6, -14, -24, -14, 10, -14, 0, 3, 5, -24, -2, -30, 3, 7, -8, 25, 17, -31, 12, -6, 7, -3, -6, -13, 8, -6, -36, -11, 41, -9, -10, -3, -27, -2, 4, -5, 1, -19, 7, -33, -9, -4, 4, -28, 10, 3, 10, 18, -16, -7, -14, 9, 23, -43, -11, 0, 8, -5, -12, -13, 0, 6, -10, 22, 11, -27, 3, 3, 2, -23, 4, 8, -10, -11, -18, 17, 22, 15, -19, 11, -22, 17, 2, 8, -12, 8, -6, -37, -19, -14, 4, -28, -3, -22, -1, 23, -10, -2, -6, 15, 21, -20, -11, 14, -7, 3, -17, -5, -9, -4, 3, -11, 1, -16, 5, 11, 6, -18, 2, 18, -6, 8, 1, -11, 18, -17, -10, 8, 6, 11, -8, 0, -4, -4, -17, -36, -20, 0, -12, -13, 8, -32, 11, 26, 4, 7, 18, 10, 10, -11, 2, -1, -20, -5, 1, -1, 0, 0, 12, 5, 2, 6, 17, 9, -8, -2, 2, 21, -7, -7, 0, -24, 14, -6, -5, -1, 4, -8, -15, -8, 4, 9, -15, 11, -4, -3, 18, -5, -2, -1, 9, 7, 6, -5, -34, -15, 15, 13, -4, 19, 2, -9, 9, -18, -2, 31, -1, 12, 0, -37, 3, 20, 16, 9, -15, -5, 5, -16, -20, -3, 35, 6, 7, 0, -17, 2, -5, 19, 14, -7, 7, 16, 7, -5, 0, -8, 0, 8, 14, 9, -11, -32, -24, 21, 16, -6, -11, 15, 7, -26, -11, -14, -4, 11, -4, 5, 13, 2, 4, 6, -2, -7, 5, 6, 7, -18, -20, 7, 27, 13, -11, 1, -27, 4, 0, -2, 6, -6, -11, -22, -13, -1, 12, -5, 5, -19, 2, 3, -9, -15, 19, 18, 12, -5, -30, -2, 9, -5, -9, -5, -13, -18, 0, 2, 4, 4, 8, 16, 2, -3, -1, 7, 13, 7, 1, -39, 30, -6, 3, -2, 14, 13, -11, -9, -8, -8, -20, -4, -2, -9, -13, -5, 16, -12, -1, 16, 3, 10, 11, 10, 6, 9, -8, 8, -31, 6, -29, -5, -3, -15, 4, 16, -5, -1, 1, -2, 6, 14, 6, 13, -10, -10, -3, 3, 2, -25, 6, 13, -5, 6, -9, -12, 1, 2, -13, 32, 20, -8, 8)
  );
  ----------------
END PACKAGE CNN_Data_Package;
